module top ;
reg [7:0] a ;
reg [7:0] b ;
 
wire [15:0] product ;
 
wallace  wa_1 (a,b,product);


initial
begin

a = 8'd0; b = 8'd0;  #10 
a = 8'd0; b = 8'd1;  #10 
a = 8'd0; b = 8'd2;  #10 
a = 8'd0; b = 8'd3;  #10 
a = 8'd0; b = 8'd4;  #10 
a = 8'd0; b = 8'd5;  #10 
a = 8'd0; b = 8'd6;  #10 
a = 8'd0; b = 8'd7;  #10 
a = 8'd0; b = 8'd8;  #10 
a = 8'd0; b = 8'd9;  #10 
a = 8'd0; b = 8'd10;  #10 
a = 8'd0; b = 8'd11;  #10 
a = 8'd0; b = 8'd12;  #10 
a = 8'd0; b = 8'd13;  #10 
a = 8'd0; b = 8'd14;  #10 
a = 8'd0; b = 8'd15;  #10 
a = 8'd0; b = 8'd16;  #10 
a = 8'd0; b = 8'd17;  #10 
a = 8'd0; b = 8'd18;  #10 
a = 8'd0; b = 8'd19;  #10 
a = 8'd0; b = 8'd20;  #10 
a = 8'd0; b = 8'd21;  #10 
a = 8'd0; b = 8'd22;  #10 
a = 8'd0; b = 8'd23;  #10 
a = 8'd0; b = 8'd24;  #10 
a = 8'd0; b = 8'd25;  #10 
a = 8'd0; b = 8'd26;  #10 
a = 8'd0; b = 8'd27;  #10 
a = 8'd0; b = 8'd28;  #10 
a = 8'd0; b = 8'd29;  #10 
a = 8'd0; b = 8'd30;  #10 
a = 8'd0; b = 8'd31;  #10 
a = 8'd0; b = 8'd32;  #10 
a = 8'd0; b = 8'd33;  #10 
a = 8'd0; b = 8'd34;  #10 
a = 8'd0; b = 8'd35;  #10 
a = 8'd0; b = 8'd36;  #10 
a = 8'd0; b = 8'd37;  #10 
a = 8'd0; b = 8'd38;  #10 
a = 8'd0; b = 8'd39;  #10 
a = 8'd0; b = 8'd40;  #10 
a = 8'd0; b = 8'd41;  #10 
a = 8'd0; b = 8'd42;  #10 
a = 8'd0; b = 8'd43;  #10 
a = 8'd0; b = 8'd44;  #10 
a = 8'd0; b = 8'd45;  #10 
a = 8'd0; b = 8'd46;  #10 
a = 8'd0; b = 8'd47;  #10 
a = 8'd0; b = 8'd48;  #10 
a = 8'd0; b = 8'd49;  #10 
a = 8'd0; b = 8'd50;  #10 
a = 8'd0; b = 8'd51;  #10 
a = 8'd0; b = 8'd52;  #10 
a = 8'd0; b = 8'd53;  #10 
a = 8'd0; b = 8'd54;  #10 
a = 8'd0; b = 8'd55;  #10 
a = 8'd0; b = 8'd56;  #10 
a = 8'd0; b = 8'd57;  #10 
a = 8'd0; b = 8'd58;  #10 
a = 8'd0; b = 8'd59;  #10 
a = 8'd0; b = 8'd60;  #10 
a = 8'd0; b = 8'd61;  #10 
a = 8'd0; b = 8'd62;  #10 
a = 8'd0; b = 8'd63;  #10 
a = 8'd0; b = 8'd64;  #10 
a = 8'd0; b = 8'd65;  #10 
a = 8'd0; b = 8'd66;  #10 
a = 8'd0; b = 8'd67;  #10 
a = 8'd0; b = 8'd68;  #10 
a = 8'd0; b = 8'd69;  #10 
a = 8'd0; b = 8'd70;  #10 
a = 8'd0; b = 8'd71;  #10 
a = 8'd0; b = 8'd72;  #10 
a = 8'd0; b = 8'd73;  #10 
a = 8'd0; b = 8'd74;  #10 
a = 8'd0; b = 8'd75;  #10 
a = 8'd0; b = 8'd76;  #10 
a = 8'd0; b = 8'd77;  #10 
a = 8'd0; b = 8'd78;  #10 
a = 8'd0; b = 8'd79;  #10 
a = 8'd0; b = 8'd80;  #10 
a = 8'd0; b = 8'd81;  #10 
a = 8'd0; b = 8'd82;  #10 
a = 8'd0; b = 8'd83;  #10 
a = 8'd0; b = 8'd84;  #10 
a = 8'd0; b = 8'd85;  #10 
a = 8'd0; b = 8'd86;  #10 
a = 8'd0; b = 8'd87;  #10 
a = 8'd0; b = 8'd88;  #10 
a = 8'd0; b = 8'd89;  #10 
a = 8'd0; b = 8'd90;  #10 
a = 8'd0; b = 8'd91;  #10 
a = 8'd0; b = 8'd92;  #10 
a = 8'd0; b = 8'd93;  #10 
a = 8'd0; b = 8'd94;  #10 
a = 8'd0; b = 8'd95;  #10 
a = 8'd0; b = 8'd96;  #10 
a = 8'd0; b = 8'd97;  #10 
a = 8'd0; b = 8'd98;  #10 
a = 8'd0; b = 8'd99;  #10 
a = 8'd0; b = 8'd100;  #10 
a = 8'd0; b = 8'd101;  #10 
a = 8'd0; b = 8'd102;  #10 
a = 8'd0; b = 8'd103;  #10 
a = 8'd0; b = 8'd104;  #10 
a = 8'd0; b = 8'd105;  #10 
a = 8'd0; b = 8'd106;  #10 
a = 8'd0; b = 8'd107;  #10 
a = 8'd0; b = 8'd108;  #10 
a = 8'd0; b = 8'd109;  #10 
a = 8'd0; b = 8'd110;  #10 
a = 8'd0; b = 8'd111;  #10 
a = 8'd0; b = 8'd112;  #10 
a = 8'd0; b = 8'd113;  #10 
a = 8'd0; b = 8'd114;  #10 
a = 8'd0; b = 8'd115;  #10 
a = 8'd0; b = 8'd116;  #10 
a = 8'd0; b = 8'd117;  #10 
a = 8'd0; b = 8'd118;  #10 
a = 8'd0; b = 8'd119;  #10 
a = 8'd0; b = 8'd120;  #10 
a = 8'd0; b = 8'd121;  #10 
a = 8'd0; b = 8'd122;  #10 
a = 8'd0; b = 8'd123;  #10 
a = 8'd0; b = 8'd124;  #10 
a = 8'd0; b = 8'd125;  #10 
a = 8'd0; b = 8'd126;  #10 
a = 8'd0; b = 8'd127;  #10 
a = 8'd0; b = 8'd128;  #10 
a = 8'd0; b = 8'd129;  #10 
a = 8'd0; b = 8'd130;  #10 
a = 8'd0; b = 8'd131;  #10 
a = 8'd0; b = 8'd132;  #10 
a = 8'd0; b = 8'd133;  #10 
a = 8'd0; b = 8'd134;  #10 
a = 8'd0; b = 8'd135;  #10 
a = 8'd0; b = 8'd136;  #10 
a = 8'd0; b = 8'd137;  #10 
a = 8'd0; b = 8'd138;  #10 
a = 8'd0; b = 8'd139;  #10 
a = 8'd0; b = 8'd140;  #10 
a = 8'd0; b = 8'd141;  #10 
a = 8'd0; b = 8'd142;  #10 
a = 8'd0; b = 8'd143;  #10 
a = 8'd0; b = 8'd144;  #10 
a = 8'd0; b = 8'd145;  #10 
a = 8'd0; b = 8'd146;  #10 
a = 8'd0; b = 8'd147;  #10 
a = 8'd0; b = 8'd148;  #10 
a = 8'd0; b = 8'd149;  #10 
a = 8'd0; b = 8'd150;  #10 
a = 8'd0; b = 8'd151;  #10 
a = 8'd0; b = 8'd152;  #10 
a = 8'd0; b = 8'd153;  #10 
a = 8'd0; b = 8'd154;  #10 
a = 8'd0; b = 8'd155;  #10 
a = 8'd0; b = 8'd156;  #10 
a = 8'd0; b = 8'd157;  #10 
a = 8'd0; b = 8'd158;  #10 
a = 8'd0; b = 8'd159;  #10 
a = 8'd0; b = 8'd160;  #10 
a = 8'd0; b = 8'd161;  #10 
a = 8'd0; b = 8'd162;  #10 
a = 8'd0; b = 8'd163;  #10 
a = 8'd0; b = 8'd164;  #10 
a = 8'd0; b = 8'd165;  #10 
a = 8'd0; b = 8'd166;  #10 
a = 8'd0; b = 8'd167;  #10 
a = 8'd0; b = 8'd168;  #10 
a = 8'd0; b = 8'd169;  #10 
a = 8'd0; b = 8'd170;  #10 
a = 8'd0; b = 8'd171;  #10 
a = 8'd0; b = 8'd172;  #10 
a = 8'd0; b = 8'd173;  #10 
a = 8'd0; b = 8'd174;  #10 
a = 8'd0; b = 8'd175;  #10 
a = 8'd0; b = 8'd176;  #10 
a = 8'd0; b = 8'd177;  #10 
a = 8'd0; b = 8'd178;  #10 
a = 8'd0; b = 8'd179;  #10 
a = 8'd0; b = 8'd180;  #10 
a = 8'd0; b = 8'd181;  #10 
a = 8'd0; b = 8'd182;  #10 
a = 8'd0; b = 8'd183;  #10 
a = 8'd0; b = 8'd184;  #10 
a = 8'd0; b = 8'd185;  #10 
a = 8'd0; b = 8'd186;  #10 
a = 8'd0; b = 8'd187;  #10 
a = 8'd0; b = 8'd188;  #10 
a = 8'd0; b = 8'd189;  #10 
a = 8'd0; b = 8'd190;  #10 
a = 8'd0; b = 8'd191;  #10 
a = 8'd0; b = 8'd192;  #10 
a = 8'd0; b = 8'd193;  #10 
a = 8'd0; b = 8'd194;  #10 
a = 8'd0; b = 8'd195;  #10 
a = 8'd0; b = 8'd196;  #10 
a = 8'd0; b = 8'd197;  #10 
a = 8'd0; b = 8'd198;  #10 
a = 8'd0; b = 8'd199;  #10 
a = 8'd0; b = 8'd200;  #10 
a = 8'd0; b = 8'd201;  #10 
a = 8'd0; b = 8'd202;  #10 
a = 8'd0; b = 8'd203;  #10 
a = 8'd0; b = 8'd204;  #10 
a = 8'd0; b = 8'd205;  #10 
a = 8'd0; b = 8'd206;  #10 
a = 8'd0; b = 8'd207;  #10 
a = 8'd0; b = 8'd208;  #10 
a = 8'd0; b = 8'd209;  #10 
a = 8'd0; b = 8'd210;  #10 
a = 8'd0; b = 8'd211;  #10 
a = 8'd0; b = 8'd212;  #10 
a = 8'd0; b = 8'd213;  #10 
a = 8'd0; b = 8'd214;  #10 
a = 8'd0; b = 8'd215;  #10 
a = 8'd0; b = 8'd216;  #10 
a = 8'd0; b = 8'd217;  #10 
a = 8'd0; b = 8'd218;  #10 
a = 8'd0; b = 8'd219;  #10 
a = 8'd0; b = 8'd220;  #10 
a = 8'd0; b = 8'd221;  #10 
a = 8'd0; b = 8'd222;  #10 
a = 8'd0; b = 8'd223;  #10 
a = 8'd0; b = 8'd224;  #10 
a = 8'd0; b = 8'd225;  #10 
a = 8'd0; b = 8'd226;  #10 
a = 8'd0; b = 8'd227;  #10 
a = 8'd0; b = 8'd228;  #10 
a = 8'd0; b = 8'd229;  #10 
a = 8'd0; b = 8'd230;  #10 
a = 8'd0; b = 8'd231;  #10 
a = 8'd0; b = 8'd232;  #10 
a = 8'd0; b = 8'd233;  #10 
a = 8'd0; b = 8'd234;  #10 
a = 8'd0; b = 8'd235;  #10 
a = 8'd0; b = 8'd236;  #10 
a = 8'd0; b = 8'd237;  #10 
a = 8'd0; b = 8'd238;  #10 
a = 8'd0; b = 8'd239;  #10 
a = 8'd0; b = 8'd240;  #10 
a = 8'd0; b = 8'd241;  #10 
a = 8'd0; b = 8'd242;  #10 
a = 8'd0; b = 8'd243;  #10 
a = 8'd0; b = 8'd244;  #10 
a = 8'd0; b = 8'd245;  #10 
a = 8'd0; b = 8'd246;  #10 
a = 8'd0; b = 8'd247;  #10 
a = 8'd0; b = 8'd248;  #10 
a = 8'd0; b = 8'd249;  #10 
a = 8'd0; b = 8'd250;  #10 
a = 8'd0; b = 8'd251;  #10 
a = 8'd0; b = 8'd252;  #10 
a = 8'd0; b = 8'd253;  #10 
a = 8'd0; b = 8'd254;  #10 
a = 8'd0; b = 8'd255;  #10 
a = 8'd1; b = 8'd0;  #10 
a = 8'd1; b = 8'd1;  #10 
a = 8'd1; b = 8'd2;  #10 
a = 8'd1; b = 8'd3;  #10 
a = 8'd1; b = 8'd4;  #10 
a = 8'd1; b = 8'd5;  #10 
a = 8'd1; b = 8'd6;  #10 
a = 8'd1; b = 8'd7;  #10 
a = 8'd1; b = 8'd8;  #10 
a = 8'd1; b = 8'd9;  #10 
a = 8'd1; b = 8'd10;  #10 
a = 8'd1; b = 8'd11;  #10 
a = 8'd1; b = 8'd12;  #10 
a = 8'd1; b = 8'd13;  #10 
a = 8'd1; b = 8'd14;  #10 
a = 8'd1; b = 8'd15;  #10 
a = 8'd1; b = 8'd16;  #10 
a = 8'd1; b = 8'd17;  #10 
a = 8'd1; b = 8'd18;  #10 
a = 8'd1; b = 8'd19;  #10 
a = 8'd1; b = 8'd20;  #10 
a = 8'd1; b = 8'd21;  #10 
a = 8'd1; b = 8'd22;  #10 
a = 8'd1; b = 8'd23;  #10 
a = 8'd1; b = 8'd24;  #10 
a = 8'd1; b = 8'd25;  #10 
a = 8'd1; b = 8'd26;  #10 
a = 8'd1; b = 8'd27;  #10 
a = 8'd1; b = 8'd28;  #10 
a = 8'd1; b = 8'd29;  #10 
a = 8'd1; b = 8'd30;  #10 
a = 8'd1; b = 8'd31;  #10 
a = 8'd1; b = 8'd32;  #10 
a = 8'd1; b = 8'd33;  #10 
a = 8'd1; b = 8'd34;  #10 
a = 8'd1; b = 8'd35;  #10 
a = 8'd1; b = 8'd36;  #10 
a = 8'd1; b = 8'd37;  #10 
a = 8'd1; b = 8'd38;  #10 
a = 8'd1; b = 8'd39;  #10 
a = 8'd1; b = 8'd40;  #10 
a = 8'd1; b = 8'd41;  #10 
a = 8'd1; b = 8'd42;  #10 
a = 8'd1; b = 8'd43;  #10 
a = 8'd1; b = 8'd44;  #10 
a = 8'd1; b = 8'd45;  #10 
a = 8'd1; b = 8'd46;  #10 
a = 8'd1; b = 8'd47;  #10 
a = 8'd1; b = 8'd48;  #10 
a = 8'd1; b = 8'd49;  #10 
a = 8'd1; b = 8'd50;  #10 
a = 8'd1; b = 8'd51;  #10 
a = 8'd1; b = 8'd52;  #10 
a = 8'd1; b = 8'd53;  #10 
a = 8'd1; b = 8'd54;  #10 
a = 8'd1; b = 8'd55;  #10 
a = 8'd1; b = 8'd56;  #10 
a = 8'd1; b = 8'd57;  #10 
a = 8'd1; b = 8'd58;  #10 
a = 8'd1; b = 8'd59;  #10 
a = 8'd1; b = 8'd60;  #10 
a = 8'd1; b = 8'd61;  #10 
a = 8'd1; b = 8'd62;  #10 
a = 8'd1; b = 8'd63;  #10 
a = 8'd1; b = 8'd64;  #10 
a = 8'd1; b = 8'd65;  #10 
a = 8'd1; b = 8'd66;  #10 
a = 8'd1; b = 8'd67;  #10 
a = 8'd1; b = 8'd68;  #10 
a = 8'd1; b = 8'd69;  #10 
a = 8'd1; b = 8'd70;  #10 
a = 8'd1; b = 8'd71;  #10 
a = 8'd1; b = 8'd72;  #10 
a = 8'd1; b = 8'd73;  #10 
a = 8'd1; b = 8'd74;  #10 
a = 8'd1; b = 8'd75;  #10 
a = 8'd1; b = 8'd76;  #10 
a = 8'd1; b = 8'd77;  #10 
a = 8'd1; b = 8'd78;  #10 
a = 8'd1; b = 8'd79;  #10 
a = 8'd1; b = 8'd80;  #10 
a = 8'd1; b = 8'd81;  #10 
a = 8'd1; b = 8'd82;  #10 
a = 8'd1; b = 8'd83;  #10 
a = 8'd1; b = 8'd84;  #10 
a = 8'd1; b = 8'd85;  #10 
a = 8'd1; b = 8'd86;  #10 
a = 8'd1; b = 8'd87;  #10 
a = 8'd1; b = 8'd88;  #10 
a = 8'd1; b = 8'd89;  #10 
a = 8'd1; b = 8'd90;  #10 
a = 8'd1; b = 8'd91;  #10 
a = 8'd1; b = 8'd92;  #10 
a = 8'd1; b = 8'd93;  #10 
a = 8'd1; b = 8'd94;  #10 
a = 8'd1; b = 8'd95;  #10 
a = 8'd1; b = 8'd96;  #10 
a = 8'd1; b = 8'd97;  #10 
a = 8'd1; b = 8'd98;  #10 
a = 8'd1; b = 8'd99;  #10 
a = 8'd1; b = 8'd100;  #10 
a = 8'd1; b = 8'd101;  #10 
a = 8'd1; b = 8'd102;  #10 
a = 8'd1; b = 8'd103;  #10 
a = 8'd1; b = 8'd104;  #10 
a = 8'd1; b = 8'd105;  #10 
a = 8'd1; b = 8'd106;  #10 
a = 8'd1; b = 8'd107;  #10 
a = 8'd1; b = 8'd108;  #10 
a = 8'd1; b = 8'd109;  #10 
a = 8'd1; b = 8'd110;  #10 
a = 8'd1; b = 8'd111;  #10 
a = 8'd1; b = 8'd112;  #10 
a = 8'd1; b = 8'd113;  #10 
a = 8'd1; b = 8'd114;  #10 
a = 8'd1; b = 8'd115;  #10 
a = 8'd1; b = 8'd116;  #10 
a = 8'd1; b = 8'd117;  #10 
a = 8'd1; b = 8'd118;  #10 
a = 8'd1; b = 8'd119;  #10 
a = 8'd1; b = 8'd120;  #10 
a = 8'd1; b = 8'd121;  #10 
a = 8'd1; b = 8'd122;  #10 
a = 8'd1; b = 8'd123;  #10 
a = 8'd1; b = 8'd124;  #10 
a = 8'd1; b = 8'd125;  #10 
a = 8'd1; b = 8'd126;  #10 
a = 8'd1; b = 8'd127;  #10 
a = 8'd1; b = 8'd128;  #10 
a = 8'd1; b = 8'd129;  #10 
a = 8'd1; b = 8'd130;  #10 
a = 8'd1; b = 8'd131;  #10 
a = 8'd1; b = 8'd132;  #10 
a = 8'd1; b = 8'd133;  #10 
a = 8'd1; b = 8'd134;  #10 
a = 8'd1; b = 8'd135;  #10 
a = 8'd1; b = 8'd136;  #10 
a = 8'd1; b = 8'd137;  #10 
a = 8'd1; b = 8'd138;  #10 
a = 8'd1; b = 8'd139;  #10 
a = 8'd1; b = 8'd140;  #10 
a = 8'd1; b = 8'd141;  #10 
a = 8'd1; b = 8'd142;  #10 
a = 8'd1; b = 8'd143;  #10 
a = 8'd1; b = 8'd144;  #10 
a = 8'd1; b = 8'd145;  #10 
a = 8'd1; b = 8'd146;  #10 
a = 8'd1; b = 8'd147;  #10 
a = 8'd1; b = 8'd148;  #10 
a = 8'd1; b = 8'd149;  #10 
a = 8'd1; b = 8'd150;  #10 
a = 8'd1; b = 8'd151;  #10 
a = 8'd1; b = 8'd152;  #10 
a = 8'd1; b = 8'd153;  #10 
a = 8'd1; b = 8'd154;  #10 
a = 8'd1; b = 8'd155;  #10 
a = 8'd1; b = 8'd156;  #10 
a = 8'd1; b = 8'd157;  #10 
a = 8'd1; b = 8'd158;  #10 
a = 8'd1; b = 8'd159;  #10 
a = 8'd1; b = 8'd160;  #10 
a = 8'd1; b = 8'd161;  #10 
a = 8'd1; b = 8'd162;  #10 
a = 8'd1; b = 8'd163;  #10 
a = 8'd1; b = 8'd164;  #10 
a = 8'd1; b = 8'd165;  #10 
a = 8'd1; b = 8'd166;  #10 
a = 8'd1; b = 8'd167;  #10 
a = 8'd1; b = 8'd168;  #10 
a = 8'd1; b = 8'd169;  #10 
a = 8'd1; b = 8'd170;  #10 
a = 8'd1; b = 8'd171;  #10 
a = 8'd1; b = 8'd172;  #10 
a = 8'd1; b = 8'd173;  #10 
a = 8'd1; b = 8'd174;  #10 
a = 8'd1; b = 8'd175;  #10 
a = 8'd1; b = 8'd176;  #10 
a = 8'd1; b = 8'd177;  #10 
a = 8'd1; b = 8'd178;  #10 
a = 8'd1; b = 8'd179;  #10 
a = 8'd1; b = 8'd180;  #10 
a = 8'd1; b = 8'd181;  #10 
a = 8'd1; b = 8'd182;  #10 
a = 8'd1; b = 8'd183;  #10 
a = 8'd1; b = 8'd184;  #10 
a = 8'd1; b = 8'd185;  #10 
a = 8'd1; b = 8'd186;  #10 
a = 8'd1; b = 8'd187;  #10 
a = 8'd1; b = 8'd188;  #10 
a = 8'd1; b = 8'd189;  #10 
a = 8'd1; b = 8'd190;  #10 
a = 8'd1; b = 8'd191;  #10 
a = 8'd1; b = 8'd192;  #10 
a = 8'd1; b = 8'd193;  #10 
a = 8'd1; b = 8'd194;  #10 
a = 8'd1; b = 8'd195;  #10 
a = 8'd1; b = 8'd196;  #10 
a = 8'd1; b = 8'd197;  #10 
a = 8'd1; b = 8'd198;  #10 
a = 8'd1; b = 8'd199;  #10 
a = 8'd1; b = 8'd200;  #10 
a = 8'd1; b = 8'd201;  #10 
a = 8'd1; b = 8'd202;  #10 
a = 8'd1; b = 8'd203;  #10 
a = 8'd1; b = 8'd204;  #10 
a = 8'd1; b = 8'd205;  #10 
a = 8'd1; b = 8'd206;  #10 
a = 8'd1; b = 8'd207;  #10 
a = 8'd1; b = 8'd208;  #10 
a = 8'd1; b = 8'd209;  #10 
a = 8'd1; b = 8'd210;  #10 
a = 8'd1; b = 8'd211;  #10 
a = 8'd1; b = 8'd212;  #10 
a = 8'd1; b = 8'd213;  #10 
a = 8'd1; b = 8'd214;  #10 
a = 8'd1; b = 8'd215;  #10 
a = 8'd1; b = 8'd216;  #10 
a = 8'd1; b = 8'd217;  #10 
a = 8'd1; b = 8'd218;  #10 
a = 8'd1; b = 8'd219;  #10 
a = 8'd1; b = 8'd220;  #10 
a = 8'd1; b = 8'd221;  #10 
a = 8'd1; b = 8'd222;  #10 
a = 8'd1; b = 8'd223;  #10 
a = 8'd1; b = 8'd224;  #10 
a = 8'd1; b = 8'd225;  #10 
a = 8'd1; b = 8'd226;  #10 
a = 8'd1; b = 8'd227;  #10 
a = 8'd1; b = 8'd228;  #10 
a = 8'd1; b = 8'd229;  #10 
a = 8'd1; b = 8'd230;  #10 
a = 8'd1; b = 8'd231;  #10 
a = 8'd1; b = 8'd232;  #10 
a = 8'd1; b = 8'd233;  #10 
a = 8'd1; b = 8'd234;  #10 
a = 8'd1; b = 8'd235;  #10 
a = 8'd1; b = 8'd236;  #10 
a = 8'd1; b = 8'd237;  #10 
a = 8'd1; b = 8'd238;  #10 
a = 8'd1; b = 8'd239;  #10 
a = 8'd1; b = 8'd240;  #10 
a = 8'd1; b = 8'd241;  #10 
a = 8'd1; b = 8'd242;  #10 
a = 8'd1; b = 8'd243;  #10 
a = 8'd1; b = 8'd244;  #10 
a = 8'd1; b = 8'd245;  #10 
a = 8'd1; b = 8'd246;  #10 
a = 8'd1; b = 8'd247;  #10 
a = 8'd1; b = 8'd248;  #10 
a = 8'd1; b = 8'd249;  #10 
a = 8'd1; b = 8'd250;  #10 
a = 8'd1; b = 8'd251;  #10 
a = 8'd1; b = 8'd252;  #10 
a = 8'd1; b = 8'd253;  #10 
a = 8'd1; b = 8'd254;  #10 
a = 8'd1; b = 8'd255;  #10 
a = 8'd2; b = 8'd0;  #10 
a = 8'd2; b = 8'd1;  #10 
a = 8'd2; b = 8'd2;  #10 
a = 8'd2; b = 8'd3;  #10 
a = 8'd2; b = 8'd4;  #10 
a = 8'd2; b = 8'd5;  #10 
a = 8'd2; b = 8'd6;  #10 
a = 8'd2; b = 8'd7;  #10 
a = 8'd2; b = 8'd8;  #10 
a = 8'd2; b = 8'd9;  #10 
a = 8'd2; b = 8'd10;  #10 
a = 8'd2; b = 8'd11;  #10 
a = 8'd2; b = 8'd12;  #10 
a = 8'd2; b = 8'd13;  #10 
a = 8'd2; b = 8'd14;  #10 
a = 8'd2; b = 8'd15;  #10 
a = 8'd2; b = 8'd16;  #10 
a = 8'd2; b = 8'd17;  #10 
a = 8'd2; b = 8'd18;  #10 
a = 8'd2; b = 8'd19;  #10 
a = 8'd2; b = 8'd20;  #10 
a = 8'd2; b = 8'd21;  #10 
a = 8'd2; b = 8'd22;  #10 
a = 8'd2; b = 8'd23;  #10 
a = 8'd2; b = 8'd24;  #10 
a = 8'd2; b = 8'd25;  #10 
a = 8'd2; b = 8'd26;  #10 
a = 8'd2; b = 8'd27;  #10 
a = 8'd2; b = 8'd28;  #10 
a = 8'd2; b = 8'd29;  #10 
a = 8'd2; b = 8'd30;  #10 
a = 8'd2; b = 8'd31;  #10 
a = 8'd2; b = 8'd32;  #10 
a = 8'd2; b = 8'd33;  #10 
a = 8'd2; b = 8'd34;  #10 
a = 8'd2; b = 8'd35;  #10 
a = 8'd2; b = 8'd36;  #10 
a = 8'd2; b = 8'd37;  #10 
a = 8'd2; b = 8'd38;  #10 
a = 8'd2; b = 8'd39;  #10 
a = 8'd2; b = 8'd40;  #10 
a = 8'd2; b = 8'd41;  #10 
a = 8'd2; b = 8'd42;  #10 
a = 8'd2; b = 8'd43;  #10 
a = 8'd2; b = 8'd44;  #10 
a = 8'd2; b = 8'd45;  #10 
a = 8'd2; b = 8'd46;  #10 
a = 8'd2; b = 8'd47;  #10 
a = 8'd2; b = 8'd48;  #10 
a = 8'd2; b = 8'd49;  #10 
a = 8'd2; b = 8'd50;  #10 
a = 8'd2; b = 8'd51;  #10 
a = 8'd2; b = 8'd52;  #10 
a = 8'd2; b = 8'd53;  #10 
a = 8'd2; b = 8'd54;  #10 
a = 8'd2; b = 8'd55;  #10 
a = 8'd2; b = 8'd56;  #10 
a = 8'd2; b = 8'd57;  #10 
a = 8'd2; b = 8'd58;  #10 
a = 8'd2; b = 8'd59;  #10 
a = 8'd2; b = 8'd60;  #10 
a = 8'd2; b = 8'd61;  #10 
a = 8'd2; b = 8'd62;  #10 
a = 8'd2; b = 8'd63;  #10 
a = 8'd2; b = 8'd64;  #10 
a = 8'd2; b = 8'd65;  #10 
a = 8'd2; b = 8'd66;  #10 
a = 8'd2; b = 8'd67;  #10 
a = 8'd2; b = 8'd68;  #10 
a = 8'd2; b = 8'd69;  #10 
a = 8'd2; b = 8'd70;  #10 
a = 8'd2; b = 8'd71;  #10 
a = 8'd2; b = 8'd72;  #10 
a = 8'd2; b = 8'd73;  #10 
a = 8'd2; b = 8'd74;  #10 
a = 8'd2; b = 8'd75;  #10 
a = 8'd2; b = 8'd76;  #10 
a = 8'd2; b = 8'd77;  #10 
a = 8'd2; b = 8'd78;  #10 
a = 8'd2; b = 8'd79;  #10 
a = 8'd2; b = 8'd80;  #10 
a = 8'd2; b = 8'd81;  #10 
a = 8'd2; b = 8'd82;  #10 
a = 8'd2; b = 8'd83;  #10 
a = 8'd2; b = 8'd84;  #10 
a = 8'd2; b = 8'd85;  #10 
a = 8'd2; b = 8'd86;  #10 
a = 8'd2; b = 8'd87;  #10 
a = 8'd2; b = 8'd88;  #10 
a = 8'd2; b = 8'd89;  #10 
a = 8'd2; b = 8'd90;  #10 
a = 8'd2; b = 8'd91;  #10 
a = 8'd2; b = 8'd92;  #10 
a = 8'd2; b = 8'd93;  #10 
a = 8'd2; b = 8'd94;  #10 
a = 8'd2; b = 8'd95;  #10 
a = 8'd2; b = 8'd96;  #10 
a = 8'd2; b = 8'd97;  #10 
a = 8'd2; b = 8'd98;  #10 
a = 8'd2; b = 8'd99;  #10 
a = 8'd2; b = 8'd100;  #10 
a = 8'd2; b = 8'd101;  #10 
a = 8'd2; b = 8'd102;  #10 
a = 8'd2; b = 8'd103;  #10 
a = 8'd2; b = 8'd104;  #10 
a = 8'd2; b = 8'd105;  #10 
a = 8'd2; b = 8'd106;  #10 
a = 8'd2; b = 8'd107;  #10 
a = 8'd2; b = 8'd108;  #10 
a = 8'd2; b = 8'd109;  #10 
a = 8'd2; b = 8'd110;  #10 
a = 8'd2; b = 8'd111;  #10 
a = 8'd2; b = 8'd112;  #10 
a = 8'd2; b = 8'd113;  #10 
a = 8'd2; b = 8'd114;  #10 
a = 8'd2; b = 8'd115;  #10 
a = 8'd2; b = 8'd116;  #10 
a = 8'd2; b = 8'd117;  #10 
a = 8'd2; b = 8'd118;  #10 
a = 8'd2; b = 8'd119;  #10 
a = 8'd2; b = 8'd120;  #10 
a = 8'd2; b = 8'd121;  #10 
a = 8'd2; b = 8'd122;  #10 
a = 8'd2; b = 8'd123;  #10 
a = 8'd2; b = 8'd124;  #10 
a = 8'd2; b = 8'd125;  #10 
a = 8'd2; b = 8'd126;  #10 
a = 8'd2; b = 8'd127;  #10 
a = 8'd2; b = 8'd128;  #10 
a = 8'd2; b = 8'd129;  #10 
a = 8'd2; b = 8'd130;  #10 
a = 8'd2; b = 8'd131;  #10 
a = 8'd2; b = 8'd132;  #10 
a = 8'd2; b = 8'd133;  #10 
a = 8'd2; b = 8'd134;  #10 
a = 8'd2; b = 8'd135;  #10 
a = 8'd2; b = 8'd136;  #10 
a = 8'd2; b = 8'd137;  #10 
a = 8'd2; b = 8'd138;  #10 
a = 8'd2; b = 8'd139;  #10 
a = 8'd2; b = 8'd140;  #10 
a = 8'd2; b = 8'd141;  #10 
a = 8'd2; b = 8'd142;  #10 
a = 8'd2; b = 8'd143;  #10 
a = 8'd2; b = 8'd144;  #10 
a = 8'd2; b = 8'd145;  #10 
a = 8'd2; b = 8'd146;  #10 
a = 8'd2; b = 8'd147;  #10 
a = 8'd2; b = 8'd148;  #10 
a = 8'd2; b = 8'd149;  #10 
a = 8'd2; b = 8'd150;  #10 
a = 8'd2; b = 8'd151;  #10 
a = 8'd2; b = 8'd152;  #10 
a = 8'd2; b = 8'd153;  #10 
a = 8'd2; b = 8'd154;  #10 
a = 8'd2; b = 8'd155;  #10 
a = 8'd2; b = 8'd156;  #10 
a = 8'd2; b = 8'd157;  #10 
a = 8'd2; b = 8'd158;  #10 
a = 8'd2; b = 8'd159;  #10 
a = 8'd2; b = 8'd160;  #10 
a = 8'd2; b = 8'd161;  #10 
a = 8'd2; b = 8'd162;  #10 
a = 8'd2; b = 8'd163;  #10 
a = 8'd2; b = 8'd164;  #10 
a = 8'd2; b = 8'd165;  #10 
a = 8'd2; b = 8'd166;  #10 
a = 8'd2; b = 8'd167;  #10 
a = 8'd2; b = 8'd168;  #10 
a = 8'd2; b = 8'd169;  #10 
a = 8'd2; b = 8'd170;  #10 
a = 8'd2; b = 8'd171;  #10 
a = 8'd2; b = 8'd172;  #10 
a = 8'd2; b = 8'd173;  #10 
a = 8'd2; b = 8'd174;  #10 
a = 8'd2; b = 8'd175;  #10 
a = 8'd2; b = 8'd176;  #10 
a = 8'd2; b = 8'd177;  #10 
a = 8'd2; b = 8'd178;  #10 
a = 8'd2; b = 8'd179;  #10 
a = 8'd2; b = 8'd180;  #10 
a = 8'd2; b = 8'd181;  #10 
a = 8'd2; b = 8'd182;  #10 
a = 8'd2; b = 8'd183;  #10 
a = 8'd2; b = 8'd184;  #10 
a = 8'd2; b = 8'd185;  #10 
a = 8'd2; b = 8'd186;  #10 
a = 8'd2; b = 8'd187;  #10 
a = 8'd2; b = 8'd188;  #10 
a = 8'd2; b = 8'd189;  #10 
a = 8'd2; b = 8'd190;  #10 
a = 8'd2; b = 8'd191;  #10 
a = 8'd2; b = 8'd192;  #10 
a = 8'd2; b = 8'd193;  #10 
a = 8'd2; b = 8'd194;  #10 
a = 8'd2; b = 8'd195;  #10 
a = 8'd2; b = 8'd196;  #10 
a = 8'd2; b = 8'd197;  #10 
a = 8'd2; b = 8'd198;  #10 
a = 8'd2; b = 8'd199;  #10 
a = 8'd2; b = 8'd200;  #10 
a = 8'd2; b = 8'd201;  #10 
a = 8'd2; b = 8'd202;  #10 
a = 8'd2; b = 8'd203;  #10 
a = 8'd2; b = 8'd204;  #10 
a = 8'd2; b = 8'd205;  #10 
a = 8'd2; b = 8'd206;  #10 
a = 8'd2; b = 8'd207;  #10 
a = 8'd2; b = 8'd208;  #10 
a = 8'd2; b = 8'd209;  #10 
a = 8'd2; b = 8'd210;  #10 
a = 8'd2; b = 8'd211;  #10 
a = 8'd2; b = 8'd212;  #10 
a = 8'd2; b = 8'd213;  #10 
a = 8'd2; b = 8'd214;  #10 
a = 8'd2; b = 8'd215;  #10 
a = 8'd2; b = 8'd216;  #10 
a = 8'd2; b = 8'd217;  #10 
a = 8'd2; b = 8'd218;  #10 
a = 8'd2; b = 8'd219;  #10 
a = 8'd2; b = 8'd220;  #10 
a = 8'd2; b = 8'd221;  #10 
a = 8'd2; b = 8'd222;  #10 
a = 8'd2; b = 8'd223;  #10 
a = 8'd2; b = 8'd224;  #10 
a = 8'd2; b = 8'd225;  #10 
a = 8'd2; b = 8'd226;  #10 
a = 8'd2; b = 8'd227;  #10 
a = 8'd2; b = 8'd228;  #10 
a = 8'd2; b = 8'd229;  #10 
a = 8'd2; b = 8'd230;  #10 
a = 8'd2; b = 8'd231;  #10 
a = 8'd2; b = 8'd232;  #10 
a = 8'd2; b = 8'd233;  #10 
a = 8'd2; b = 8'd234;  #10 
a = 8'd2; b = 8'd235;  #10 
a = 8'd2; b = 8'd236;  #10 
a = 8'd2; b = 8'd237;  #10 
a = 8'd2; b = 8'd238;  #10 
a = 8'd2; b = 8'd239;  #10 
a = 8'd2; b = 8'd240;  #10 
a = 8'd2; b = 8'd241;  #10 
a = 8'd2; b = 8'd242;  #10 
a = 8'd2; b = 8'd243;  #10 
a = 8'd2; b = 8'd244;  #10 
a = 8'd2; b = 8'd245;  #10 
a = 8'd2; b = 8'd246;  #10 
a = 8'd2; b = 8'd247;  #10 
a = 8'd2; b = 8'd248;  #10 
a = 8'd2; b = 8'd249;  #10 
a = 8'd2; b = 8'd250;  #10 
a = 8'd2; b = 8'd251;  #10 
a = 8'd2; b = 8'd252;  #10 
a = 8'd2; b = 8'd253;  #10 
a = 8'd2; b = 8'd254;  #10 
a = 8'd2; b = 8'd255;  #10 
a = 8'd3; b = 8'd0;  #10 
a = 8'd3; b = 8'd1;  #10 
a = 8'd3; b = 8'd2;  #10 
a = 8'd3; b = 8'd3;  #10 
a = 8'd3; b = 8'd4;  #10 
a = 8'd3; b = 8'd5;  #10 
a = 8'd3; b = 8'd6;  #10 
a = 8'd3; b = 8'd7;  #10 
a = 8'd3; b = 8'd8;  #10 
a = 8'd3; b = 8'd9;  #10 
a = 8'd3; b = 8'd10;  #10 
a = 8'd3; b = 8'd11;  #10 
a = 8'd3; b = 8'd12;  #10 
a = 8'd3; b = 8'd13;  #10 
a = 8'd3; b = 8'd14;  #10 
a = 8'd3; b = 8'd15;  #10 
a = 8'd3; b = 8'd16;  #10 
a = 8'd3; b = 8'd17;  #10 
a = 8'd3; b = 8'd18;  #10 
a = 8'd3; b = 8'd19;  #10 
a = 8'd3; b = 8'd20;  #10 
a = 8'd3; b = 8'd21;  #10 
a = 8'd3; b = 8'd22;  #10 
a = 8'd3; b = 8'd23;  #10 
a = 8'd3; b = 8'd24;  #10 
a = 8'd3; b = 8'd25;  #10 
a = 8'd3; b = 8'd26;  #10 
a = 8'd3; b = 8'd27;  #10 
a = 8'd3; b = 8'd28;  #10 
a = 8'd3; b = 8'd29;  #10 
a = 8'd3; b = 8'd30;  #10 
a = 8'd3; b = 8'd31;  #10 
a = 8'd3; b = 8'd32;  #10 
a = 8'd3; b = 8'd33;  #10 
a = 8'd3; b = 8'd34;  #10 
a = 8'd3; b = 8'd35;  #10 
a = 8'd3; b = 8'd36;  #10 
a = 8'd3; b = 8'd37;  #10 
a = 8'd3; b = 8'd38;  #10 
a = 8'd3; b = 8'd39;  #10 
a = 8'd3; b = 8'd40;  #10 
a = 8'd3; b = 8'd41;  #10 
a = 8'd3; b = 8'd42;  #10 
a = 8'd3; b = 8'd43;  #10 
a = 8'd3; b = 8'd44;  #10 
a = 8'd3; b = 8'd45;  #10 
a = 8'd3; b = 8'd46;  #10 
a = 8'd3; b = 8'd47;  #10 
a = 8'd3; b = 8'd48;  #10 
a = 8'd3; b = 8'd49;  #10 
a = 8'd3; b = 8'd50;  #10 
a = 8'd3; b = 8'd51;  #10 
a = 8'd3; b = 8'd52;  #10 
a = 8'd3; b = 8'd53;  #10 
a = 8'd3; b = 8'd54;  #10 
a = 8'd3; b = 8'd55;  #10 
a = 8'd3; b = 8'd56;  #10 
a = 8'd3; b = 8'd57;  #10 
a = 8'd3; b = 8'd58;  #10 
a = 8'd3; b = 8'd59;  #10 
a = 8'd3; b = 8'd60;  #10 
a = 8'd3; b = 8'd61;  #10 
a = 8'd3; b = 8'd62;  #10 
a = 8'd3; b = 8'd63;  #10 
a = 8'd3; b = 8'd64;  #10 
a = 8'd3; b = 8'd65;  #10 
a = 8'd3; b = 8'd66;  #10 
a = 8'd3; b = 8'd67;  #10 
a = 8'd3; b = 8'd68;  #10 
a = 8'd3; b = 8'd69;  #10 
a = 8'd3; b = 8'd70;  #10 
a = 8'd3; b = 8'd71;  #10 
a = 8'd3; b = 8'd72;  #10 
a = 8'd3; b = 8'd73;  #10 
a = 8'd3; b = 8'd74;  #10 
a = 8'd3; b = 8'd75;  #10 
a = 8'd3; b = 8'd76;  #10 
a = 8'd3; b = 8'd77;  #10 
a = 8'd3; b = 8'd78;  #10 
a = 8'd3; b = 8'd79;  #10 
a = 8'd3; b = 8'd80;  #10 
a = 8'd3; b = 8'd81;  #10 
a = 8'd3; b = 8'd82;  #10 
a = 8'd3; b = 8'd83;  #10 
a = 8'd3; b = 8'd84;  #10 
a = 8'd3; b = 8'd85;  #10 
a = 8'd3; b = 8'd86;  #10 
a = 8'd3; b = 8'd87;  #10 
a = 8'd3; b = 8'd88;  #10 
a = 8'd3; b = 8'd89;  #10 
a = 8'd3; b = 8'd90;  #10 
a = 8'd3; b = 8'd91;  #10 
a = 8'd3; b = 8'd92;  #10 
a = 8'd3; b = 8'd93;  #10 
a = 8'd3; b = 8'd94;  #10 
a = 8'd3; b = 8'd95;  #10 
a = 8'd3; b = 8'd96;  #10 
a = 8'd3; b = 8'd97;  #10 
a = 8'd3; b = 8'd98;  #10 
a = 8'd3; b = 8'd99;  #10 
a = 8'd3; b = 8'd100;  #10 
a = 8'd3; b = 8'd101;  #10 
a = 8'd3; b = 8'd102;  #10 
a = 8'd3; b = 8'd103;  #10 
a = 8'd3; b = 8'd104;  #10 
a = 8'd3; b = 8'd105;  #10 
a = 8'd3; b = 8'd106;  #10 
a = 8'd3; b = 8'd107;  #10 
a = 8'd3; b = 8'd108;  #10 
a = 8'd3; b = 8'd109;  #10 
a = 8'd3; b = 8'd110;  #10 
a = 8'd3; b = 8'd111;  #10 
a = 8'd3; b = 8'd112;  #10 
a = 8'd3; b = 8'd113;  #10 
a = 8'd3; b = 8'd114;  #10 
a = 8'd3; b = 8'd115;  #10 
a = 8'd3; b = 8'd116;  #10 
a = 8'd3; b = 8'd117;  #10 
a = 8'd3; b = 8'd118;  #10 
a = 8'd3; b = 8'd119;  #10 
a = 8'd3; b = 8'd120;  #10 
a = 8'd3; b = 8'd121;  #10 
a = 8'd3; b = 8'd122;  #10 
a = 8'd3; b = 8'd123;  #10 
a = 8'd3; b = 8'd124;  #10 
a = 8'd3; b = 8'd125;  #10 
a = 8'd3; b = 8'd126;  #10 
a = 8'd3; b = 8'd127;  #10 
a = 8'd3; b = 8'd128;  #10 
a = 8'd3; b = 8'd129;  #10 
a = 8'd3; b = 8'd130;  #10 
a = 8'd3; b = 8'd131;  #10 
a = 8'd3; b = 8'd132;  #10 
a = 8'd3; b = 8'd133;  #10 
a = 8'd3; b = 8'd134;  #10 
a = 8'd3; b = 8'd135;  #10 
a = 8'd3; b = 8'd136;  #10 
a = 8'd3; b = 8'd137;  #10 
a = 8'd3; b = 8'd138;  #10 
a = 8'd3; b = 8'd139;  #10 
a = 8'd3; b = 8'd140;  #10 
a = 8'd3; b = 8'd141;  #10 
a = 8'd3; b = 8'd142;  #10 
a = 8'd3; b = 8'd143;  #10 
a = 8'd3; b = 8'd144;  #10 
a = 8'd3; b = 8'd145;  #10 
a = 8'd3; b = 8'd146;  #10 
a = 8'd3; b = 8'd147;  #10 
a = 8'd3; b = 8'd148;  #10 
a = 8'd3; b = 8'd149;  #10 
a = 8'd3; b = 8'd150;  #10 
a = 8'd3; b = 8'd151;  #10 
a = 8'd3; b = 8'd152;  #10 
a = 8'd3; b = 8'd153;  #10 
a = 8'd3; b = 8'd154;  #10 
a = 8'd3; b = 8'd155;  #10 
a = 8'd3; b = 8'd156;  #10 
a = 8'd3; b = 8'd157;  #10 
a = 8'd3; b = 8'd158;  #10 
a = 8'd3; b = 8'd159;  #10 
a = 8'd3; b = 8'd160;  #10 
a = 8'd3; b = 8'd161;  #10 
a = 8'd3; b = 8'd162;  #10 
a = 8'd3; b = 8'd163;  #10 
a = 8'd3; b = 8'd164;  #10 
a = 8'd3; b = 8'd165;  #10 
a = 8'd3; b = 8'd166;  #10 
a = 8'd3; b = 8'd167;  #10 
a = 8'd3; b = 8'd168;  #10 
a = 8'd3; b = 8'd169;  #10 
a = 8'd3; b = 8'd170;  #10 
a = 8'd3; b = 8'd171;  #10 
a = 8'd3; b = 8'd172;  #10 
a = 8'd3; b = 8'd173;  #10 
a = 8'd3; b = 8'd174;  #10 
a = 8'd3; b = 8'd175;  #10 
a = 8'd3; b = 8'd176;  #10 
a = 8'd3; b = 8'd177;  #10 
a = 8'd3; b = 8'd178;  #10 
a = 8'd3; b = 8'd179;  #10 
a = 8'd3; b = 8'd180;  #10 
a = 8'd3; b = 8'd181;  #10 
a = 8'd3; b = 8'd182;  #10 
a = 8'd3; b = 8'd183;  #10 
a = 8'd3; b = 8'd184;  #10 
a = 8'd3; b = 8'd185;  #10 
a = 8'd3; b = 8'd186;  #10 
a = 8'd3; b = 8'd187;  #10 
a = 8'd3; b = 8'd188;  #10 
a = 8'd3; b = 8'd189;  #10 
a = 8'd3; b = 8'd190;  #10 
a = 8'd3; b = 8'd191;  #10 
a = 8'd3; b = 8'd192;  #10 
a = 8'd3; b = 8'd193;  #10 
a = 8'd3; b = 8'd194;  #10 
a = 8'd3; b = 8'd195;  #10 
a = 8'd3; b = 8'd196;  #10 
a = 8'd3; b = 8'd197;  #10 
a = 8'd3; b = 8'd198;  #10 
a = 8'd3; b = 8'd199;  #10 
a = 8'd3; b = 8'd200;  #10 
a = 8'd3; b = 8'd201;  #10 
a = 8'd3; b = 8'd202;  #10 
a = 8'd3; b = 8'd203;  #10 
a = 8'd3; b = 8'd204;  #10 
a = 8'd3; b = 8'd205;  #10 
a = 8'd3; b = 8'd206;  #10 
a = 8'd3; b = 8'd207;  #10 
a = 8'd3; b = 8'd208;  #10 
a = 8'd3; b = 8'd209;  #10 
a = 8'd3; b = 8'd210;  #10 
a = 8'd3; b = 8'd211;  #10 
a = 8'd3; b = 8'd212;  #10 
a = 8'd3; b = 8'd213;  #10 
a = 8'd3; b = 8'd214;  #10 
a = 8'd3; b = 8'd215;  #10 
a = 8'd3; b = 8'd216;  #10 
a = 8'd3; b = 8'd217;  #10 
a = 8'd3; b = 8'd218;  #10 
a = 8'd3; b = 8'd219;  #10 
a = 8'd3; b = 8'd220;  #10 
a = 8'd3; b = 8'd221;  #10 
a = 8'd3; b = 8'd222;  #10 
a = 8'd3; b = 8'd223;  #10 
a = 8'd3; b = 8'd224;  #10 
a = 8'd3; b = 8'd225;  #10 
a = 8'd3; b = 8'd226;  #10 
a = 8'd3; b = 8'd227;  #10 
a = 8'd3; b = 8'd228;  #10 
a = 8'd3; b = 8'd229;  #10 
a = 8'd3; b = 8'd230;  #10 
a = 8'd3; b = 8'd231;  #10 
a = 8'd3; b = 8'd232;  #10 
a = 8'd3; b = 8'd233;  #10 
a = 8'd3; b = 8'd234;  #10 
a = 8'd3; b = 8'd235;  #10 
a = 8'd3; b = 8'd236;  #10 
a = 8'd3; b = 8'd237;  #10 
a = 8'd3; b = 8'd238;  #10 
a = 8'd3; b = 8'd239;  #10 
a = 8'd3; b = 8'd240;  #10 
a = 8'd3; b = 8'd241;  #10 
a = 8'd3; b = 8'd242;  #10 
a = 8'd3; b = 8'd243;  #10 
a = 8'd3; b = 8'd244;  #10 
a = 8'd3; b = 8'd245;  #10 
a = 8'd3; b = 8'd246;  #10 
a = 8'd3; b = 8'd247;  #10 
a = 8'd3; b = 8'd248;  #10 
a = 8'd3; b = 8'd249;  #10 
a = 8'd3; b = 8'd250;  #10 
a = 8'd3; b = 8'd251;  #10 
a = 8'd3; b = 8'd252;  #10 
a = 8'd3; b = 8'd253;  #10 
a = 8'd3; b = 8'd254;  #10 
a = 8'd3; b = 8'd255;  #10 
a = 8'd4; b = 8'd0;  #10 
a = 8'd4; b = 8'd1;  #10 
a = 8'd4; b = 8'd2;  #10 
a = 8'd4; b = 8'd3;  #10 
a = 8'd4; b = 8'd4;  #10 
a = 8'd4; b = 8'd5;  #10 
a = 8'd4; b = 8'd6;  #10 
a = 8'd4; b = 8'd7;  #10 
a = 8'd4; b = 8'd8;  #10 
a = 8'd4; b = 8'd9;  #10 
a = 8'd4; b = 8'd10;  #10 
a = 8'd4; b = 8'd11;  #10 
a = 8'd4; b = 8'd12;  #10 
a = 8'd4; b = 8'd13;  #10 
a = 8'd4; b = 8'd14;  #10 
a = 8'd4; b = 8'd15;  #10 
a = 8'd4; b = 8'd16;  #10 
a = 8'd4; b = 8'd17;  #10 
a = 8'd4; b = 8'd18;  #10 
a = 8'd4; b = 8'd19;  #10 
a = 8'd4; b = 8'd20;  #10 
a = 8'd4; b = 8'd21;  #10 
a = 8'd4; b = 8'd22;  #10 
a = 8'd4; b = 8'd23;  #10 
a = 8'd4; b = 8'd24;  #10 
a = 8'd4; b = 8'd25;  #10 
a = 8'd4; b = 8'd26;  #10 
a = 8'd4; b = 8'd27;  #10 
a = 8'd4; b = 8'd28;  #10 
a = 8'd4; b = 8'd29;  #10 
a = 8'd4; b = 8'd30;  #10 
a = 8'd4; b = 8'd31;  #10 
a = 8'd4; b = 8'd32;  #10 
a = 8'd4; b = 8'd33;  #10 
a = 8'd4; b = 8'd34;  #10 
a = 8'd4; b = 8'd35;  #10 
a = 8'd4; b = 8'd36;  #10 
a = 8'd4; b = 8'd37;  #10 
a = 8'd4; b = 8'd38;  #10 
a = 8'd4; b = 8'd39;  #10 
a = 8'd4; b = 8'd40;  #10 
a = 8'd4; b = 8'd41;  #10 
a = 8'd4; b = 8'd42;  #10 
a = 8'd4; b = 8'd43;  #10 
a = 8'd4; b = 8'd44;  #10 
a = 8'd4; b = 8'd45;  #10 
a = 8'd4; b = 8'd46;  #10 
a = 8'd4; b = 8'd47;  #10 
a = 8'd4; b = 8'd48;  #10 
a = 8'd4; b = 8'd49;  #10 
a = 8'd4; b = 8'd50;  #10 
a = 8'd4; b = 8'd51;  #10 
a = 8'd4; b = 8'd52;  #10 
a = 8'd4; b = 8'd53;  #10 
a = 8'd4; b = 8'd54;  #10 
a = 8'd4; b = 8'd55;  #10 
a = 8'd4; b = 8'd56;  #10 
a = 8'd4; b = 8'd57;  #10 
a = 8'd4; b = 8'd58;  #10 
a = 8'd4; b = 8'd59;  #10 
a = 8'd4; b = 8'd60;  #10 
a = 8'd4; b = 8'd61;  #10 
a = 8'd4; b = 8'd62;  #10 
a = 8'd4; b = 8'd63;  #10 
a = 8'd4; b = 8'd64;  #10 
a = 8'd4; b = 8'd65;  #10 
a = 8'd4; b = 8'd66;  #10 
a = 8'd4; b = 8'd67;  #10 
a = 8'd4; b = 8'd68;  #10 
a = 8'd4; b = 8'd69;  #10 
a = 8'd4; b = 8'd70;  #10 
a = 8'd4; b = 8'd71;  #10 
a = 8'd4; b = 8'd72;  #10 
a = 8'd4; b = 8'd73;  #10 
a = 8'd4; b = 8'd74;  #10 
a = 8'd4; b = 8'd75;  #10 
a = 8'd4; b = 8'd76;  #10 
a = 8'd4; b = 8'd77;  #10 
a = 8'd4; b = 8'd78;  #10 
a = 8'd4; b = 8'd79;  #10 
a = 8'd4; b = 8'd80;  #10 
a = 8'd4; b = 8'd81;  #10 
a = 8'd4; b = 8'd82;  #10 
a = 8'd4; b = 8'd83;  #10 
a = 8'd4; b = 8'd84;  #10 
a = 8'd4; b = 8'd85;  #10 
a = 8'd4; b = 8'd86;  #10 
a = 8'd4; b = 8'd87;  #10 
a = 8'd4; b = 8'd88;  #10 
a = 8'd4; b = 8'd89;  #10 
a = 8'd4; b = 8'd90;  #10 
a = 8'd4; b = 8'd91;  #10 
a = 8'd4; b = 8'd92;  #10 
a = 8'd4; b = 8'd93;  #10 
a = 8'd4; b = 8'd94;  #10 
a = 8'd4; b = 8'd95;  #10 
a = 8'd4; b = 8'd96;  #10 
a = 8'd4; b = 8'd97;  #10 
a = 8'd4; b = 8'd98;  #10 
a = 8'd4; b = 8'd99;  #10 
a = 8'd4; b = 8'd100;  #10 
a = 8'd4; b = 8'd101;  #10 
a = 8'd4; b = 8'd102;  #10 
a = 8'd4; b = 8'd103;  #10 
a = 8'd4; b = 8'd104;  #10 
a = 8'd4; b = 8'd105;  #10 
a = 8'd4; b = 8'd106;  #10 
a = 8'd4; b = 8'd107;  #10 
a = 8'd4; b = 8'd108;  #10 
a = 8'd4; b = 8'd109;  #10 
a = 8'd4; b = 8'd110;  #10 
a = 8'd4; b = 8'd111;  #10 
a = 8'd4; b = 8'd112;  #10 
a = 8'd4; b = 8'd113;  #10 
a = 8'd4; b = 8'd114;  #10 
a = 8'd4; b = 8'd115;  #10 
a = 8'd4; b = 8'd116;  #10 
a = 8'd4; b = 8'd117;  #10 
a = 8'd4; b = 8'd118;  #10 
a = 8'd4; b = 8'd119;  #10 
a = 8'd4; b = 8'd120;  #10 
a = 8'd4; b = 8'd121;  #10 
a = 8'd4; b = 8'd122;  #10 
a = 8'd4; b = 8'd123;  #10 
a = 8'd4; b = 8'd124;  #10 
a = 8'd4; b = 8'd125;  #10 
a = 8'd4; b = 8'd126;  #10 
a = 8'd4; b = 8'd127;  #10 
a = 8'd4; b = 8'd128;  #10 
a = 8'd4; b = 8'd129;  #10 
a = 8'd4; b = 8'd130;  #10 
a = 8'd4; b = 8'd131;  #10 
a = 8'd4; b = 8'd132;  #10 
a = 8'd4; b = 8'd133;  #10 
a = 8'd4; b = 8'd134;  #10 
a = 8'd4; b = 8'd135;  #10 
a = 8'd4; b = 8'd136;  #10 
a = 8'd4; b = 8'd137;  #10 
a = 8'd4; b = 8'd138;  #10 
a = 8'd4; b = 8'd139;  #10 
a = 8'd4; b = 8'd140;  #10 
a = 8'd4; b = 8'd141;  #10 
a = 8'd4; b = 8'd142;  #10 
a = 8'd4; b = 8'd143;  #10 
a = 8'd4; b = 8'd144;  #10 
a = 8'd4; b = 8'd145;  #10 
a = 8'd4; b = 8'd146;  #10 
a = 8'd4; b = 8'd147;  #10 
a = 8'd4; b = 8'd148;  #10 
a = 8'd4; b = 8'd149;  #10 
a = 8'd4; b = 8'd150;  #10 
a = 8'd4; b = 8'd151;  #10 
a = 8'd4; b = 8'd152;  #10 
a = 8'd4; b = 8'd153;  #10 
a = 8'd4; b = 8'd154;  #10 
a = 8'd4; b = 8'd155;  #10 
a = 8'd4; b = 8'd156;  #10 
a = 8'd4; b = 8'd157;  #10 
a = 8'd4; b = 8'd158;  #10 
a = 8'd4; b = 8'd159;  #10 
a = 8'd4; b = 8'd160;  #10 
a = 8'd4; b = 8'd161;  #10 
a = 8'd4; b = 8'd162;  #10 
a = 8'd4; b = 8'd163;  #10 
a = 8'd4; b = 8'd164;  #10 
a = 8'd4; b = 8'd165;  #10 
a = 8'd4; b = 8'd166;  #10 
a = 8'd4; b = 8'd167;  #10 
a = 8'd4; b = 8'd168;  #10 
a = 8'd4; b = 8'd169;  #10 
a = 8'd4; b = 8'd170;  #10 
a = 8'd4; b = 8'd171;  #10 
a = 8'd4; b = 8'd172;  #10 
a = 8'd4; b = 8'd173;  #10 
a = 8'd4; b = 8'd174;  #10 
a = 8'd4; b = 8'd175;  #10 
a = 8'd4; b = 8'd176;  #10 
a = 8'd4; b = 8'd177;  #10 
a = 8'd4; b = 8'd178;  #10 
a = 8'd4; b = 8'd179;  #10 
a = 8'd4; b = 8'd180;  #10 
a = 8'd4; b = 8'd181;  #10 
a = 8'd4; b = 8'd182;  #10 
a = 8'd4; b = 8'd183;  #10 
a = 8'd4; b = 8'd184;  #10 
a = 8'd4; b = 8'd185;  #10 
a = 8'd4; b = 8'd186;  #10 
a = 8'd4; b = 8'd187;  #10 
a = 8'd4; b = 8'd188;  #10 
a = 8'd4; b = 8'd189;  #10 
a = 8'd4; b = 8'd190;  #10 
a = 8'd4; b = 8'd191;  #10 
a = 8'd4; b = 8'd192;  #10 
a = 8'd4; b = 8'd193;  #10 
a = 8'd4; b = 8'd194;  #10 
a = 8'd4; b = 8'd195;  #10 
a = 8'd4; b = 8'd196;  #10 
a = 8'd4; b = 8'd197;  #10 
a = 8'd4; b = 8'd198;  #10 
a = 8'd4; b = 8'd199;  #10 
a = 8'd4; b = 8'd200;  #10 
a = 8'd4; b = 8'd201;  #10 
a = 8'd4; b = 8'd202;  #10 
a = 8'd4; b = 8'd203;  #10 
a = 8'd4; b = 8'd204;  #10 
a = 8'd4; b = 8'd205;  #10 
a = 8'd4; b = 8'd206;  #10 
a = 8'd4; b = 8'd207;  #10 
a = 8'd4; b = 8'd208;  #10 
a = 8'd4; b = 8'd209;  #10 
a = 8'd4; b = 8'd210;  #10 
a = 8'd4; b = 8'd211;  #10 
a = 8'd4; b = 8'd212;  #10 
a = 8'd4; b = 8'd213;  #10 
a = 8'd4; b = 8'd214;  #10 
a = 8'd4; b = 8'd215;  #10 
a = 8'd4; b = 8'd216;  #10 
a = 8'd4; b = 8'd217;  #10 
a = 8'd4; b = 8'd218;  #10 
a = 8'd4; b = 8'd219;  #10 
a = 8'd4; b = 8'd220;  #10 
a = 8'd4; b = 8'd221;  #10 
a = 8'd4; b = 8'd222;  #10 
a = 8'd4; b = 8'd223;  #10 
a = 8'd4; b = 8'd224;  #10 
a = 8'd4; b = 8'd225;  #10 
a = 8'd4; b = 8'd226;  #10 
a = 8'd4; b = 8'd227;  #10 
a = 8'd4; b = 8'd228;  #10 
a = 8'd4; b = 8'd229;  #10 
a = 8'd4; b = 8'd230;  #10 
a = 8'd4; b = 8'd231;  #10 
a = 8'd4; b = 8'd232;  #10 
a = 8'd4; b = 8'd233;  #10 
a = 8'd4; b = 8'd234;  #10 
a = 8'd4; b = 8'd235;  #10 
a = 8'd4; b = 8'd236;  #10 
a = 8'd4; b = 8'd237;  #10 
a = 8'd4; b = 8'd238;  #10 
a = 8'd4; b = 8'd239;  #10 
a = 8'd4; b = 8'd240;  #10 
a = 8'd4; b = 8'd241;  #10 
a = 8'd4; b = 8'd242;  #10 
a = 8'd4; b = 8'd243;  #10 
a = 8'd4; b = 8'd244;  #10 
a = 8'd4; b = 8'd245;  #10 
a = 8'd4; b = 8'd246;  #10 
a = 8'd4; b = 8'd247;  #10 
a = 8'd4; b = 8'd248;  #10 
a = 8'd4; b = 8'd249;  #10 
a = 8'd4; b = 8'd250;  #10 
a = 8'd4; b = 8'd251;  #10 
a = 8'd4; b = 8'd252;  #10 
a = 8'd4; b = 8'd253;  #10 
a = 8'd4; b = 8'd254;  #10 
a = 8'd4; b = 8'd255;  #10 
a = 8'd5; b = 8'd0;  #10 
a = 8'd5; b = 8'd1;  #10 
a = 8'd5; b = 8'd2;  #10 
a = 8'd5; b = 8'd3;  #10 
a = 8'd5; b = 8'd4;  #10 
a = 8'd5; b = 8'd5;  #10 
a = 8'd5; b = 8'd6;  #10 
a = 8'd5; b = 8'd7;  #10 
a = 8'd5; b = 8'd8;  #10 
a = 8'd5; b = 8'd9;  #10 
a = 8'd5; b = 8'd10;  #10 
a = 8'd5; b = 8'd11;  #10 
a = 8'd5; b = 8'd12;  #10 
a = 8'd5; b = 8'd13;  #10 
a = 8'd5; b = 8'd14;  #10 
a = 8'd5; b = 8'd15;  #10 
a = 8'd5; b = 8'd16;  #10 
a = 8'd5; b = 8'd17;  #10 
a = 8'd5; b = 8'd18;  #10 
a = 8'd5; b = 8'd19;  #10 
a = 8'd5; b = 8'd20;  #10 
a = 8'd5; b = 8'd21;  #10 
a = 8'd5; b = 8'd22;  #10 
a = 8'd5; b = 8'd23;  #10 
a = 8'd5; b = 8'd24;  #10 
a = 8'd5; b = 8'd25;  #10 
a = 8'd5; b = 8'd26;  #10 
a = 8'd5; b = 8'd27;  #10 
a = 8'd5; b = 8'd28;  #10 
a = 8'd5; b = 8'd29;  #10 
a = 8'd5; b = 8'd30;  #10 
a = 8'd5; b = 8'd31;  #10 
a = 8'd5; b = 8'd32;  #10 
a = 8'd5; b = 8'd33;  #10 
a = 8'd5; b = 8'd34;  #10 
a = 8'd5; b = 8'd35;  #10 
a = 8'd5; b = 8'd36;  #10 
a = 8'd5; b = 8'd37;  #10 
a = 8'd5; b = 8'd38;  #10 
a = 8'd5; b = 8'd39;  #10 
a = 8'd5; b = 8'd40;  #10 
a = 8'd5; b = 8'd41;  #10 
a = 8'd5; b = 8'd42;  #10 
a = 8'd5; b = 8'd43;  #10 
a = 8'd5; b = 8'd44;  #10 
a = 8'd5; b = 8'd45;  #10 
a = 8'd5; b = 8'd46;  #10 
a = 8'd5; b = 8'd47;  #10 
a = 8'd5; b = 8'd48;  #10 
a = 8'd5; b = 8'd49;  #10 
a = 8'd5; b = 8'd50;  #10 
a = 8'd5; b = 8'd51;  #10 
a = 8'd5; b = 8'd52;  #10 
a = 8'd5; b = 8'd53;  #10 
a = 8'd5; b = 8'd54;  #10 
a = 8'd5; b = 8'd55;  #10 
a = 8'd5; b = 8'd56;  #10 
a = 8'd5; b = 8'd57;  #10 
a = 8'd5; b = 8'd58;  #10 
a = 8'd5; b = 8'd59;  #10 
a = 8'd5; b = 8'd60;  #10 
a = 8'd5; b = 8'd61;  #10 
a = 8'd5; b = 8'd62;  #10 
a = 8'd5; b = 8'd63;  #10 
a = 8'd5; b = 8'd64;  #10 
a = 8'd5; b = 8'd65;  #10 
a = 8'd5; b = 8'd66;  #10 
a = 8'd5; b = 8'd67;  #10 
a = 8'd5; b = 8'd68;  #10 
a = 8'd5; b = 8'd69;  #10 
a = 8'd5; b = 8'd70;  #10 
a = 8'd5; b = 8'd71;  #10 
a = 8'd5; b = 8'd72;  #10 
a = 8'd5; b = 8'd73;  #10 
a = 8'd5; b = 8'd74;  #10 
a = 8'd5; b = 8'd75;  #10 
a = 8'd5; b = 8'd76;  #10 
a = 8'd5; b = 8'd77;  #10 
a = 8'd5; b = 8'd78;  #10 
a = 8'd5; b = 8'd79;  #10 
a = 8'd5; b = 8'd80;  #10 
a = 8'd5; b = 8'd81;  #10 
a = 8'd5; b = 8'd82;  #10 
a = 8'd5; b = 8'd83;  #10 
a = 8'd5; b = 8'd84;  #10 
a = 8'd5; b = 8'd85;  #10 
a = 8'd5; b = 8'd86;  #10 
a = 8'd5; b = 8'd87;  #10 
a = 8'd5; b = 8'd88;  #10 
a = 8'd5; b = 8'd89;  #10 
a = 8'd5; b = 8'd90;  #10 
a = 8'd5; b = 8'd91;  #10 
a = 8'd5; b = 8'd92;  #10 
a = 8'd5; b = 8'd93;  #10 
a = 8'd5; b = 8'd94;  #10 
a = 8'd5; b = 8'd95;  #10 
a = 8'd5; b = 8'd96;  #10 
a = 8'd5; b = 8'd97;  #10 
a = 8'd5; b = 8'd98;  #10 
a = 8'd5; b = 8'd99;  #10 
a = 8'd5; b = 8'd100;  #10 
a = 8'd5; b = 8'd101;  #10 
a = 8'd5; b = 8'd102;  #10 
a = 8'd5; b = 8'd103;  #10 
a = 8'd5; b = 8'd104;  #10 
a = 8'd5; b = 8'd105;  #10 
a = 8'd5; b = 8'd106;  #10 
a = 8'd5; b = 8'd107;  #10 
a = 8'd5; b = 8'd108;  #10 
a = 8'd5; b = 8'd109;  #10 
a = 8'd5; b = 8'd110;  #10 
a = 8'd5; b = 8'd111;  #10 
a = 8'd5; b = 8'd112;  #10 
a = 8'd5; b = 8'd113;  #10 
a = 8'd5; b = 8'd114;  #10 
a = 8'd5; b = 8'd115;  #10 
a = 8'd5; b = 8'd116;  #10 
a = 8'd5; b = 8'd117;  #10 
a = 8'd5; b = 8'd118;  #10 
a = 8'd5; b = 8'd119;  #10 
a = 8'd5; b = 8'd120;  #10 
a = 8'd5; b = 8'd121;  #10 
a = 8'd5; b = 8'd122;  #10 
a = 8'd5; b = 8'd123;  #10 
a = 8'd5; b = 8'd124;  #10 
a = 8'd5; b = 8'd125;  #10 
a = 8'd5; b = 8'd126;  #10 
a = 8'd5; b = 8'd127;  #10 
a = 8'd5; b = 8'd128;  #10 
a = 8'd5; b = 8'd129;  #10 
a = 8'd5; b = 8'd130;  #10 
a = 8'd5; b = 8'd131;  #10 
a = 8'd5; b = 8'd132;  #10 
a = 8'd5; b = 8'd133;  #10 
a = 8'd5; b = 8'd134;  #10 
a = 8'd5; b = 8'd135;  #10 
a = 8'd5; b = 8'd136;  #10 
a = 8'd5; b = 8'd137;  #10 
a = 8'd5; b = 8'd138;  #10 
a = 8'd5; b = 8'd139;  #10 
a = 8'd5; b = 8'd140;  #10 
a = 8'd5; b = 8'd141;  #10 
a = 8'd5; b = 8'd142;  #10 
a = 8'd5; b = 8'd143;  #10 
a = 8'd5; b = 8'd144;  #10 
a = 8'd5; b = 8'd145;  #10 
a = 8'd5; b = 8'd146;  #10 
a = 8'd5; b = 8'd147;  #10 
a = 8'd5; b = 8'd148;  #10 
a = 8'd5; b = 8'd149;  #10 
a = 8'd5; b = 8'd150;  #10 
a = 8'd5; b = 8'd151;  #10 
a = 8'd5; b = 8'd152;  #10 
a = 8'd5; b = 8'd153;  #10 
a = 8'd5; b = 8'd154;  #10 
a = 8'd5; b = 8'd155;  #10 
a = 8'd5; b = 8'd156;  #10 
a = 8'd5; b = 8'd157;  #10 
a = 8'd5; b = 8'd158;  #10 
a = 8'd5; b = 8'd159;  #10 
a = 8'd5; b = 8'd160;  #10 
a = 8'd5; b = 8'd161;  #10 
a = 8'd5; b = 8'd162;  #10 
a = 8'd5; b = 8'd163;  #10 
a = 8'd5; b = 8'd164;  #10 
a = 8'd5; b = 8'd165;  #10 
a = 8'd5; b = 8'd166;  #10 
a = 8'd5; b = 8'd167;  #10 
a = 8'd5; b = 8'd168;  #10 
a = 8'd5; b = 8'd169;  #10 
a = 8'd5; b = 8'd170;  #10 
a = 8'd5; b = 8'd171;  #10 
a = 8'd5; b = 8'd172;  #10 
a = 8'd5; b = 8'd173;  #10 
a = 8'd5; b = 8'd174;  #10 
a = 8'd5; b = 8'd175;  #10 
a = 8'd5; b = 8'd176;  #10 
a = 8'd5; b = 8'd177;  #10 
a = 8'd5; b = 8'd178;  #10 
a = 8'd5; b = 8'd179;  #10 
a = 8'd5; b = 8'd180;  #10 
a = 8'd5; b = 8'd181;  #10 
a = 8'd5; b = 8'd182;  #10 
a = 8'd5; b = 8'd183;  #10 
a = 8'd5; b = 8'd184;  #10 
a = 8'd5; b = 8'd185;  #10 
a = 8'd5; b = 8'd186;  #10 
a = 8'd5; b = 8'd187;  #10 
a = 8'd5; b = 8'd188;  #10 
a = 8'd5; b = 8'd189;  #10 
a = 8'd5; b = 8'd190;  #10 
a = 8'd5; b = 8'd191;  #10 
a = 8'd5; b = 8'd192;  #10 
a = 8'd5; b = 8'd193;  #10 
a = 8'd5; b = 8'd194;  #10 
a = 8'd5; b = 8'd195;  #10 
a = 8'd5; b = 8'd196;  #10 
a = 8'd5; b = 8'd197;  #10 
a = 8'd5; b = 8'd198;  #10 
a = 8'd5; b = 8'd199;  #10 
a = 8'd5; b = 8'd200;  #10 
a = 8'd5; b = 8'd201;  #10 
a = 8'd5; b = 8'd202;  #10 
a = 8'd5; b = 8'd203;  #10 
a = 8'd5; b = 8'd204;  #10 
a = 8'd5; b = 8'd205;  #10 
a = 8'd5; b = 8'd206;  #10 
a = 8'd5; b = 8'd207;  #10 
a = 8'd5; b = 8'd208;  #10 
a = 8'd5; b = 8'd209;  #10 
a = 8'd5; b = 8'd210;  #10 
a = 8'd5; b = 8'd211;  #10 
a = 8'd5; b = 8'd212;  #10 
a = 8'd5; b = 8'd213;  #10 
a = 8'd5; b = 8'd214;  #10 
a = 8'd5; b = 8'd215;  #10 
a = 8'd5; b = 8'd216;  #10 
a = 8'd5; b = 8'd217;  #10 
a = 8'd5; b = 8'd218;  #10 
a = 8'd5; b = 8'd219;  #10 
a = 8'd5; b = 8'd220;  #10 
a = 8'd5; b = 8'd221;  #10 
a = 8'd5; b = 8'd222;  #10 
a = 8'd5; b = 8'd223;  #10 
a = 8'd5; b = 8'd224;  #10 
a = 8'd5; b = 8'd225;  #10 
a = 8'd5; b = 8'd226;  #10 
a = 8'd5; b = 8'd227;  #10 
a = 8'd5; b = 8'd228;  #10 
a = 8'd5; b = 8'd229;  #10 
a = 8'd5; b = 8'd230;  #10 
a = 8'd5; b = 8'd231;  #10 
a = 8'd5; b = 8'd232;  #10 
a = 8'd5; b = 8'd233;  #10 
a = 8'd5; b = 8'd234;  #10 
a = 8'd5; b = 8'd235;  #10 
a = 8'd5; b = 8'd236;  #10 
a = 8'd5; b = 8'd237;  #10 
a = 8'd5; b = 8'd238;  #10 
a = 8'd5; b = 8'd239;  #10 
a = 8'd5; b = 8'd240;  #10 
a = 8'd5; b = 8'd241;  #10 
a = 8'd5; b = 8'd242;  #10 
a = 8'd5; b = 8'd243;  #10 
a = 8'd5; b = 8'd244;  #10 
a = 8'd5; b = 8'd245;  #10 
a = 8'd5; b = 8'd246;  #10 
a = 8'd5; b = 8'd247;  #10 
a = 8'd5; b = 8'd248;  #10 
a = 8'd5; b = 8'd249;  #10 
a = 8'd5; b = 8'd250;  #10 
a = 8'd5; b = 8'd251;  #10 
a = 8'd5; b = 8'd252;  #10 
a = 8'd5; b = 8'd253;  #10 
a = 8'd5; b = 8'd254;  #10 
a = 8'd5; b = 8'd255;  #10 
a = 8'd6; b = 8'd0;  #10 
a = 8'd6; b = 8'd1;  #10 
a = 8'd6; b = 8'd2;  #10 
a = 8'd6; b = 8'd3;  #10 
a = 8'd6; b = 8'd4;  #10 
a = 8'd6; b = 8'd5;  #10 
a = 8'd6; b = 8'd6;  #10 
a = 8'd6; b = 8'd7;  #10 
a = 8'd6; b = 8'd8;  #10 
a = 8'd6; b = 8'd9;  #10 
a = 8'd6; b = 8'd10;  #10 
a = 8'd6; b = 8'd11;  #10 
a = 8'd6; b = 8'd12;  #10 
a = 8'd6; b = 8'd13;  #10 
a = 8'd6; b = 8'd14;  #10 
a = 8'd6; b = 8'd15;  #10 
a = 8'd6; b = 8'd16;  #10 
a = 8'd6; b = 8'd17;  #10 
a = 8'd6; b = 8'd18;  #10 
a = 8'd6; b = 8'd19;  #10 
a = 8'd6; b = 8'd20;  #10 
a = 8'd6; b = 8'd21;  #10 
a = 8'd6; b = 8'd22;  #10 
a = 8'd6; b = 8'd23;  #10 
a = 8'd6; b = 8'd24;  #10 
a = 8'd6; b = 8'd25;  #10 
a = 8'd6; b = 8'd26;  #10 
a = 8'd6; b = 8'd27;  #10 
a = 8'd6; b = 8'd28;  #10 
a = 8'd6; b = 8'd29;  #10 
a = 8'd6; b = 8'd30;  #10 
a = 8'd6; b = 8'd31;  #10 
a = 8'd6; b = 8'd32;  #10 
a = 8'd6; b = 8'd33;  #10 
a = 8'd6; b = 8'd34;  #10 
a = 8'd6; b = 8'd35;  #10 
a = 8'd6; b = 8'd36;  #10 
a = 8'd6; b = 8'd37;  #10 
a = 8'd6; b = 8'd38;  #10 
a = 8'd6; b = 8'd39;  #10 
a = 8'd6; b = 8'd40;  #10 
a = 8'd6; b = 8'd41;  #10 
a = 8'd6; b = 8'd42;  #10 
a = 8'd6; b = 8'd43;  #10 
a = 8'd6; b = 8'd44;  #10 
a = 8'd6; b = 8'd45;  #10 
a = 8'd6; b = 8'd46;  #10 
a = 8'd6; b = 8'd47;  #10 
a = 8'd6; b = 8'd48;  #10 
a = 8'd6; b = 8'd49;  #10 
a = 8'd6; b = 8'd50;  #10 
a = 8'd6; b = 8'd51;  #10 
a = 8'd6; b = 8'd52;  #10 
a = 8'd6; b = 8'd53;  #10 
a = 8'd6; b = 8'd54;  #10 
a = 8'd6; b = 8'd55;  #10 
a = 8'd6; b = 8'd56;  #10 
a = 8'd6; b = 8'd57;  #10 
a = 8'd6; b = 8'd58;  #10 
a = 8'd6; b = 8'd59;  #10 
a = 8'd6; b = 8'd60;  #10 
a = 8'd6; b = 8'd61;  #10 
a = 8'd6; b = 8'd62;  #10 
a = 8'd6; b = 8'd63;  #10 
a = 8'd6; b = 8'd64;  #10 
a = 8'd6; b = 8'd65;  #10 
a = 8'd6; b = 8'd66;  #10 
a = 8'd6; b = 8'd67;  #10 
a = 8'd6; b = 8'd68;  #10 
a = 8'd6; b = 8'd69;  #10 
a = 8'd6; b = 8'd70;  #10 
a = 8'd6; b = 8'd71;  #10 
a = 8'd6; b = 8'd72;  #10 
a = 8'd6; b = 8'd73;  #10 
a = 8'd6; b = 8'd74;  #10 
a = 8'd6; b = 8'd75;  #10 
a = 8'd6; b = 8'd76;  #10 
a = 8'd6; b = 8'd77;  #10 
a = 8'd6; b = 8'd78;  #10 
a = 8'd6; b = 8'd79;  #10 
a = 8'd6; b = 8'd80;  #10 
a = 8'd6; b = 8'd81;  #10 
a = 8'd6; b = 8'd82;  #10 
a = 8'd6; b = 8'd83;  #10 
a = 8'd6; b = 8'd84;  #10 
a = 8'd6; b = 8'd85;  #10 
a = 8'd6; b = 8'd86;  #10 
a = 8'd6; b = 8'd87;  #10 
a = 8'd6; b = 8'd88;  #10 
a = 8'd6; b = 8'd89;  #10 
a = 8'd6; b = 8'd90;  #10 
a = 8'd6; b = 8'd91;  #10 
a = 8'd6; b = 8'd92;  #10 
a = 8'd6; b = 8'd93;  #10 
a = 8'd6; b = 8'd94;  #10 
a = 8'd6; b = 8'd95;  #10 
a = 8'd6; b = 8'd96;  #10 
a = 8'd6; b = 8'd97;  #10 
a = 8'd6; b = 8'd98;  #10 
a = 8'd6; b = 8'd99;  #10 
a = 8'd6; b = 8'd100;  #10 
a = 8'd6; b = 8'd101;  #10 
a = 8'd6; b = 8'd102;  #10 
a = 8'd6; b = 8'd103;  #10 
a = 8'd6; b = 8'd104;  #10 
a = 8'd6; b = 8'd105;  #10 
a = 8'd6; b = 8'd106;  #10 
a = 8'd6; b = 8'd107;  #10 
a = 8'd6; b = 8'd108;  #10 
a = 8'd6; b = 8'd109;  #10 
a = 8'd6; b = 8'd110;  #10 
a = 8'd6; b = 8'd111;  #10 
a = 8'd6; b = 8'd112;  #10 
a = 8'd6; b = 8'd113;  #10 
a = 8'd6; b = 8'd114;  #10 
a = 8'd6; b = 8'd115;  #10 
a = 8'd6; b = 8'd116;  #10 
a = 8'd6; b = 8'd117;  #10 
a = 8'd6; b = 8'd118;  #10 
a = 8'd6; b = 8'd119;  #10 
a = 8'd6; b = 8'd120;  #10 
a = 8'd6; b = 8'd121;  #10 
a = 8'd6; b = 8'd122;  #10 
a = 8'd6; b = 8'd123;  #10 
a = 8'd6; b = 8'd124;  #10 
a = 8'd6; b = 8'd125;  #10 
a = 8'd6; b = 8'd126;  #10 
a = 8'd6; b = 8'd127;  #10 
a = 8'd6; b = 8'd128;  #10 
a = 8'd6; b = 8'd129;  #10 
a = 8'd6; b = 8'd130;  #10 
a = 8'd6; b = 8'd131;  #10 
a = 8'd6; b = 8'd132;  #10 
a = 8'd6; b = 8'd133;  #10 
a = 8'd6; b = 8'd134;  #10 
a = 8'd6; b = 8'd135;  #10 
a = 8'd6; b = 8'd136;  #10 
a = 8'd6; b = 8'd137;  #10 
a = 8'd6; b = 8'd138;  #10 
a = 8'd6; b = 8'd139;  #10 
a = 8'd6; b = 8'd140;  #10 
a = 8'd6; b = 8'd141;  #10 
a = 8'd6; b = 8'd142;  #10 
a = 8'd6; b = 8'd143;  #10 
a = 8'd6; b = 8'd144;  #10 
a = 8'd6; b = 8'd145;  #10 
a = 8'd6; b = 8'd146;  #10 
a = 8'd6; b = 8'd147;  #10 
a = 8'd6; b = 8'd148;  #10 
a = 8'd6; b = 8'd149;  #10 
a = 8'd6; b = 8'd150;  #10 
a = 8'd6; b = 8'd151;  #10 
a = 8'd6; b = 8'd152;  #10 
a = 8'd6; b = 8'd153;  #10 
a = 8'd6; b = 8'd154;  #10 
a = 8'd6; b = 8'd155;  #10 
a = 8'd6; b = 8'd156;  #10 
a = 8'd6; b = 8'd157;  #10 
a = 8'd6; b = 8'd158;  #10 
a = 8'd6; b = 8'd159;  #10 
a = 8'd6; b = 8'd160;  #10 
a = 8'd6; b = 8'd161;  #10 
a = 8'd6; b = 8'd162;  #10 
a = 8'd6; b = 8'd163;  #10 
a = 8'd6; b = 8'd164;  #10 
a = 8'd6; b = 8'd165;  #10 
a = 8'd6; b = 8'd166;  #10 
a = 8'd6; b = 8'd167;  #10 
a = 8'd6; b = 8'd168;  #10 
a = 8'd6; b = 8'd169;  #10 
a = 8'd6; b = 8'd170;  #10 
a = 8'd6; b = 8'd171;  #10 
a = 8'd6; b = 8'd172;  #10 
a = 8'd6; b = 8'd173;  #10 
a = 8'd6; b = 8'd174;  #10 
a = 8'd6; b = 8'd175;  #10 
a = 8'd6; b = 8'd176;  #10 
a = 8'd6; b = 8'd177;  #10 
a = 8'd6; b = 8'd178;  #10 
a = 8'd6; b = 8'd179;  #10 
a = 8'd6; b = 8'd180;  #10 
a = 8'd6; b = 8'd181;  #10 
a = 8'd6; b = 8'd182;  #10 
a = 8'd6; b = 8'd183;  #10 
a = 8'd6; b = 8'd184;  #10 
a = 8'd6; b = 8'd185;  #10 
a = 8'd6; b = 8'd186;  #10 
a = 8'd6; b = 8'd187;  #10 
a = 8'd6; b = 8'd188;  #10 
a = 8'd6; b = 8'd189;  #10 
a = 8'd6; b = 8'd190;  #10 
a = 8'd6; b = 8'd191;  #10 
a = 8'd6; b = 8'd192;  #10 
a = 8'd6; b = 8'd193;  #10 
a = 8'd6; b = 8'd194;  #10 
a = 8'd6; b = 8'd195;  #10 
a = 8'd6; b = 8'd196;  #10 
a = 8'd6; b = 8'd197;  #10 
a = 8'd6; b = 8'd198;  #10 
a = 8'd6; b = 8'd199;  #10 
a = 8'd6; b = 8'd200;  #10 
a = 8'd6; b = 8'd201;  #10 
a = 8'd6; b = 8'd202;  #10 
a = 8'd6; b = 8'd203;  #10 
a = 8'd6; b = 8'd204;  #10 
a = 8'd6; b = 8'd205;  #10 
a = 8'd6; b = 8'd206;  #10 
a = 8'd6; b = 8'd207;  #10 
a = 8'd6; b = 8'd208;  #10 
a = 8'd6; b = 8'd209;  #10 
a = 8'd6; b = 8'd210;  #10 
a = 8'd6; b = 8'd211;  #10 
a = 8'd6; b = 8'd212;  #10 
a = 8'd6; b = 8'd213;  #10 
a = 8'd6; b = 8'd214;  #10 
a = 8'd6; b = 8'd215;  #10 
a = 8'd6; b = 8'd216;  #10 
a = 8'd6; b = 8'd217;  #10 
a = 8'd6; b = 8'd218;  #10 
a = 8'd6; b = 8'd219;  #10 
a = 8'd6; b = 8'd220;  #10 
a = 8'd6; b = 8'd221;  #10 
a = 8'd6; b = 8'd222;  #10 
a = 8'd6; b = 8'd223;  #10 
a = 8'd6; b = 8'd224;  #10 
a = 8'd6; b = 8'd225;  #10 
a = 8'd6; b = 8'd226;  #10 
a = 8'd6; b = 8'd227;  #10 
a = 8'd6; b = 8'd228;  #10 
a = 8'd6; b = 8'd229;  #10 
a = 8'd6; b = 8'd230;  #10 
a = 8'd6; b = 8'd231;  #10 
a = 8'd6; b = 8'd232;  #10 
a = 8'd6; b = 8'd233;  #10 
a = 8'd6; b = 8'd234;  #10 
a = 8'd6; b = 8'd235;  #10 
a = 8'd6; b = 8'd236;  #10 
a = 8'd6; b = 8'd237;  #10 
a = 8'd6; b = 8'd238;  #10 
a = 8'd6; b = 8'd239;  #10 
a = 8'd6; b = 8'd240;  #10 
a = 8'd6; b = 8'd241;  #10 
a = 8'd6; b = 8'd242;  #10 
a = 8'd6; b = 8'd243;  #10 
a = 8'd6; b = 8'd244;  #10 
a = 8'd6; b = 8'd245;  #10 
a = 8'd6; b = 8'd246;  #10 
a = 8'd6; b = 8'd247;  #10 
a = 8'd6; b = 8'd248;  #10 
a = 8'd6; b = 8'd249;  #10 
a = 8'd6; b = 8'd250;  #10 
a = 8'd6; b = 8'd251;  #10 
a = 8'd6; b = 8'd252;  #10 
a = 8'd6; b = 8'd253;  #10 
a = 8'd6; b = 8'd254;  #10 
a = 8'd6; b = 8'd255;  #10 
a = 8'd7; b = 8'd0;  #10 
a = 8'd7; b = 8'd1;  #10 
a = 8'd7; b = 8'd2;  #10 
a = 8'd7; b = 8'd3;  #10 
a = 8'd7; b = 8'd4;  #10 
a = 8'd7; b = 8'd5;  #10 
a = 8'd7; b = 8'd6;  #10 
a = 8'd7; b = 8'd7;  #10 
a = 8'd7; b = 8'd8;  #10 
a = 8'd7; b = 8'd9;  #10 
a = 8'd7; b = 8'd10;  #10 
a = 8'd7; b = 8'd11;  #10 
a = 8'd7; b = 8'd12;  #10 
a = 8'd7; b = 8'd13;  #10 
a = 8'd7; b = 8'd14;  #10 
a = 8'd7; b = 8'd15;  #10 
a = 8'd7; b = 8'd16;  #10 
a = 8'd7; b = 8'd17;  #10 
a = 8'd7; b = 8'd18;  #10 
a = 8'd7; b = 8'd19;  #10 
a = 8'd7; b = 8'd20;  #10 
a = 8'd7; b = 8'd21;  #10 
a = 8'd7; b = 8'd22;  #10 
a = 8'd7; b = 8'd23;  #10 
a = 8'd7; b = 8'd24;  #10 
a = 8'd7; b = 8'd25;  #10 
a = 8'd7; b = 8'd26;  #10 
a = 8'd7; b = 8'd27;  #10 
a = 8'd7; b = 8'd28;  #10 
a = 8'd7; b = 8'd29;  #10 
a = 8'd7; b = 8'd30;  #10 
a = 8'd7; b = 8'd31;  #10 
a = 8'd7; b = 8'd32;  #10 
a = 8'd7; b = 8'd33;  #10 
a = 8'd7; b = 8'd34;  #10 
a = 8'd7; b = 8'd35;  #10 
a = 8'd7; b = 8'd36;  #10 
a = 8'd7; b = 8'd37;  #10 
a = 8'd7; b = 8'd38;  #10 
a = 8'd7; b = 8'd39;  #10 
a = 8'd7; b = 8'd40;  #10 
a = 8'd7; b = 8'd41;  #10 
a = 8'd7; b = 8'd42;  #10 
a = 8'd7; b = 8'd43;  #10 
a = 8'd7; b = 8'd44;  #10 
a = 8'd7; b = 8'd45;  #10 
a = 8'd7; b = 8'd46;  #10 
a = 8'd7; b = 8'd47;  #10 
a = 8'd7; b = 8'd48;  #10 
a = 8'd7; b = 8'd49;  #10 
a = 8'd7; b = 8'd50;  #10 
a = 8'd7; b = 8'd51;  #10 
a = 8'd7; b = 8'd52;  #10 
a = 8'd7; b = 8'd53;  #10 
a = 8'd7; b = 8'd54;  #10 
a = 8'd7; b = 8'd55;  #10 
a = 8'd7; b = 8'd56;  #10 
a = 8'd7; b = 8'd57;  #10 
a = 8'd7; b = 8'd58;  #10 
a = 8'd7; b = 8'd59;  #10 
a = 8'd7; b = 8'd60;  #10 
a = 8'd7; b = 8'd61;  #10 
a = 8'd7; b = 8'd62;  #10 
a = 8'd7; b = 8'd63;  #10 
a = 8'd7; b = 8'd64;  #10 
a = 8'd7; b = 8'd65;  #10 
a = 8'd7; b = 8'd66;  #10 
a = 8'd7; b = 8'd67;  #10 
a = 8'd7; b = 8'd68;  #10 
a = 8'd7; b = 8'd69;  #10 
a = 8'd7; b = 8'd70;  #10 
a = 8'd7; b = 8'd71;  #10 
a = 8'd7; b = 8'd72;  #10 
a = 8'd7; b = 8'd73;  #10 
a = 8'd7; b = 8'd74;  #10 
a = 8'd7; b = 8'd75;  #10 
a = 8'd7; b = 8'd76;  #10 
a = 8'd7; b = 8'd77;  #10 
a = 8'd7; b = 8'd78;  #10 
a = 8'd7; b = 8'd79;  #10 
a = 8'd7; b = 8'd80;  #10 
a = 8'd7; b = 8'd81;  #10 
a = 8'd7; b = 8'd82;  #10 
a = 8'd7; b = 8'd83;  #10 
a = 8'd7; b = 8'd84;  #10 
a = 8'd7; b = 8'd85;  #10 
a = 8'd7; b = 8'd86;  #10 
a = 8'd7; b = 8'd87;  #10 
a = 8'd7; b = 8'd88;  #10 
a = 8'd7; b = 8'd89;  #10 
a = 8'd7; b = 8'd90;  #10 
a = 8'd7; b = 8'd91;  #10 
a = 8'd7; b = 8'd92;  #10 
a = 8'd7; b = 8'd93;  #10 
a = 8'd7; b = 8'd94;  #10 
a = 8'd7; b = 8'd95;  #10 
a = 8'd7; b = 8'd96;  #10 
a = 8'd7; b = 8'd97;  #10 
a = 8'd7; b = 8'd98;  #10 
a = 8'd7; b = 8'd99;  #10 
a = 8'd7; b = 8'd100;  #10 
a = 8'd7; b = 8'd101;  #10 
a = 8'd7; b = 8'd102;  #10 
a = 8'd7; b = 8'd103;  #10 
a = 8'd7; b = 8'd104;  #10 
a = 8'd7; b = 8'd105;  #10 
a = 8'd7; b = 8'd106;  #10 
a = 8'd7; b = 8'd107;  #10 
a = 8'd7; b = 8'd108;  #10 
a = 8'd7; b = 8'd109;  #10 
a = 8'd7; b = 8'd110;  #10 
a = 8'd7; b = 8'd111;  #10 
a = 8'd7; b = 8'd112;  #10 
a = 8'd7; b = 8'd113;  #10 
a = 8'd7; b = 8'd114;  #10 
a = 8'd7; b = 8'd115;  #10 
a = 8'd7; b = 8'd116;  #10 
a = 8'd7; b = 8'd117;  #10 
a = 8'd7; b = 8'd118;  #10 
a = 8'd7; b = 8'd119;  #10 
a = 8'd7; b = 8'd120;  #10 
a = 8'd7; b = 8'd121;  #10 
a = 8'd7; b = 8'd122;  #10 
a = 8'd7; b = 8'd123;  #10 
a = 8'd7; b = 8'd124;  #10 
a = 8'd7; b = 8'd125;  #10 
a = 8'd7; b = 8'd126;  #10 
a = 8'd7; b = 8'd127;  #10 
a = 8'd7; b = 8'd128;  #10 
a = 8'd7; b = 8'd129;  #10 
a = 8'd7; b = 8'd130;  #10 
a = 8'd7; b = 8'd131;  #10 
a = 8'd7; b = 8'd132;  #10 
a = 8'd7; b = 8'd133;  #10 
a = 8'd7; b = 8'd134;  #10 
a = 8'd7; b = 8'd135;  #10 
a = 8'd7; b = 8'd136;  #10 
a = 8'd7; b = 8'd137;  #10 
a = 8'd7; b = 8'd138;  #10 
a = 8'd7; b = 8'd139;  #10 
a = 8'd7; b = 8'd140;  #10 
a = 8'd7; b = 8'd141;  #10 
a = 8'd7; b = 8'd142;  #10 
a = 8'd7; b = 8'd143;  #10 
a = 8'd7; b = 8'd144;  #10 
a = 8'd7; b = 8'd145;  #10 
a = 8'd7; b = 8'd146;  #10 
a = 8'd7; b = 8'd147;  #10 
a = 8'd7; b = 8'd148;  #10 
a = 8'd7; b = 8'd149;  #10 
a = 8'd7; b = 8'd150;  #10 
a = 8'd7; b = 8'd151;  #10 
a = 8'd7; b = 8'd152;  #10 
a = 8'd7; b = 8'd153;  #10 
a = 8'd7; b = 8'd154;  #10 
a = 8'd7; b = 8'd155;  #10 
a = 8'd7; b = 8'd156;  #10 
a = 8'd7; b = 8'd157;  #10 
a = 8'd7; b = 8'd158;  #10 
a = 8'd7; b = 8'd159;  #10 
a = 8'd7; b = 8'd160;  #10 
a = 8'd7; b = 8'd161;  #10 
a = 8'd7; b = 8'd162;  #10 
a = 8'd7; b = 8'd163;  #10 
a = 8'd7; b = 8'd164;  #10 
a = 8'd7; b = 8'd165;  #10 
a = 8'd7; b = 8'd166;  #10 
a = 8'd7; b = 8'd167;  #10 
a = 8'd7; b = 8'd168;  #10 
a = 8'd7; b = 8'd169;  #10 
a = 8'd7; b = 8'd170;  #10 
a = 8'd7; b = 8'd171;  #10 
a = 8'd7; b = 8'd172;  #10 
a = 8'd7; b = 8'd173;  #10 
a = 8'd7; b = 8'd174;  #10 
a = 8'd7; b = 8'd175;  #10 
a = 8'd7; b = 8'd176;  #10 
a = 8'd7; b = 8'd177;  #10 
a = 8'd7; b = 8'd178;  #10 
a = 8'd7; b = 8'd179;  #10 
a = 8'd7; b = 8'd180;  #10 
a = 8'd7; b = 8'd181;  #10 
a = 8'd7; b = 8'd182;  #10 
a = 8'd7; b = 8'd183;  #10 
a = 8'd7; b = 8'd184;  #10 
a = 8'd7; b = 8'd185;  #10 
a = 8'd7; b = 8'd186;  #10 
a = 8'd7; b = 8'd187;  #10 
a = 8'd7; b = 8'd188;  #10 
a = 8'd7; b = 8'd189;  #10 
a = 8'd7; b = 8'd190;  #10 
a = 8'd7; b = 8'd191;  #10 
a = 8'd7; b = 8'd192;  #10 
a = 8'd7; b = 8'd193;  #10 
a = 8'd7; b = 8'd194;  #10 
a = 8'd7; b = 8'd195;  #10 
a = 8'd7; b = 8'd196;  #10 
a = 8'd7; b = 8'd197;  #10 
a = 8'd7; b = 8'd198;  #10 
a = 8'd7; b = 8'd199;  #10 
a = 8'd7; b = 8'd200;  #10 
a = 8'd7; b = 8'd201;  #10 
a = 8'd7; b = 8'd202;  #10 
a = 8'd7; b = 8'd203;  #10 
a = 8'd7; b = 8'd204;  #10 
a = 8'd7; b = 8'd205;  #10 
a = 8'd7; b = 8'd206;  #10 
a = 8'd7; b = 8'd207;  #10 
a = 8'd7; b = 8'd208;  #10 
a = 8'd7; b = 8'd209;  #10 
a = 8'd7; b = 8'd210;  #10 
a = 8'd7; b = 8'd211;  #10 
a = 8'd7; b = 8'd212;  #10 
a = 8'd7; b = 8'd213;  #10 
a = 8'd7; b = 8'd214;  #10 
a = 8'd7; b = 8'd215;  #10 
a = 8'd7; b = 8'd216;  #10 
a = 8'd7; b = 8'd217;  #10 
a = 8'd7; b = 8'd218;  #10 
a = 8'd7; b = 8'd219;  #10 
a = 8'd7; b = 8'd220;  #10 
a = 8'd7; b = 8'd221;  #10 
a = 8'd7; b = 8'd222;  #10 
a = 8'd7; b = 8'd223;  #10 
a = 8'd7; b = 8'd224;  #10 
a = 8'd7; b = 8'd225;  #10 
a = 8'd7; b = 8'd226;  #10 
a = 8'd7; b = 8'd227;  #10 
a = 8'd7; b = 8'd228;  #10 
a = 8'd7; b = 8'd229;  #10 
a = 8'd7; b = 8'd230;  #10 
a = 8'd7; b = 8'd231;  #10 
a = 8'd7; b = 8'd232;  #10 
a = 8'd7; b = 8'd233;  #10 
a = 8'd7; b = 8'd234;  #10 
a = 8'd7; b = 8'd235;  #10 
a = 8'd7; b = 8'd236;  #10 
a = 8'd7; b = 8'd237;  #10 
a = 8'd7; b = 8'd238;  #10 
a = 8'd7; b = 8'd239;  #10 
a = 8'd7; b = 8'd240;  #10 
a = 8'd7; b = 8'd241;  #10 
a = 8'd7; b = 8'd242;  #10 
a = 8'd7; b = 8'd243;  #10 
a = 8'd7; b = 8'd244;  #10 
a = 8'd7; b = 8'd245;  #10 
a = 8'd7; b = 8'd246;  #10 
a = 8'd7; b = 8'd247;  #10 
a = 8'd7; b = 8'd248;  #10 
a = 8'd7; b = 8'd249;  #10 
a = 8'd7; b = 8'd250;  #10 
a = 8'd7; b = 8'd251;  #10 
a = 8'd7; b = 8'd252;  #10 
a = 8'd7; b = 8'd253;  #10 
a = 8'd7; b = 8'd254;  #10 
a = 8'd7; b = 8'd255;  #10 
a = 8'd8; b = 8'd0;  #10 
a = 8'd8; b = 8'd1;  #10 
a = 8'd8; b = 8'd2;  #10 
a = 8'd8; b = 8'd3;  #10 
a = 8'd8; b = 8'd4;  #10 
a = 8'd8; b = 8'd5;  #10 
a = 8'd8; b = 8'd6;  #10 
a = 8'd8; b = 8'd7;  #10 
a = 8'd8; b = 8'd8;  #10 
a = 8'd8; b = 8'd9;  #10 
a = 8'd8; b = 8'd10;  #10 
a = 8'd8; b = 8'd11;  #10 
a = 8'd8; b = 8'd12;  #10 
a = 8'd8; b = 8'd13;  #10 
a = 8'd8; b = 8'd14;  #10 
a = 8'd8; b = 8'd15;  #10 
a = 8'd8; b = 8'd16;  #10 
a = 8'd8; b = 8'd17;  #10 
a = 8'd8; b = 8'd18;  #10 
a = 8'd8; b = 8'd19;  #10 
a = 8'd8; b = 8'd20;  #10 
a = 8'd8; b = 8'd21;  #10 
a = 8'd8; b = 8'd22;  #10 
a = 8'd8; b = 8'd23;  #10 
a = 8'd8; b = 8'd24;  #10 
a = 8'd8; b = 8'd25;  #10 
a = 8'd8; b = 8'd26;  #10 
a = 8'd8; b = 8'd27;  #10 
a = 8'd8; b = 8'd28;  #10 
a = 8'd8; b = 8'd29;  #10 
a = 8'd8; b = 8'd30;  #10 
a = 8'd8; b = 8'd31;  #10 
a = 8'd8; b = 8'd32;  #10 
a = 8'd8; b = 8'd33;  #10 
a = 8'd8; b = 8'd34;  #10 
a = 8'd8; b = 8'd35;  #10 
a = 8'd8; b = 8'd36;  #10 
a = 8'd8; b = 8'd37;  #10 
a = 8'd8; b = 8'd38;  #10 
a = 8'd8; b = 8'd39;  #10 
a = 8'd8; b = 8'd40;  #10 
a = 8'd8; b = 8'd41;  #10 
a = 8'd8; b = 8'd42;  #10 
a = 8'd8; b = 8'd43;  #10 
a = 8'd8; b = 8'd44;  #10 
a = 8'd8; b = 8'd45;  #10 
a = 8'd8; b = 8'd46;  #10 
a = 8'd8; b = 8'd47;  #10 
a = 8'd8; b = 8'd48;  #10 
a = 8'd8; b = 8'd49;  #10 
a = 8'd8; b = 8'd50;  #10 
a = 8'd8; b = 8'd51;  #10 
a = 8'd8; b = 8'd52;  #10 
a = 8'd8; b = 8'd53;  #10 
a = 8'd8; b = 8'd54;  #10 
a = 8'd8; b = 8'd55;  #10 
a = 8'd8; b = 8'd56;  #10 
a = 8'd8; b = 8'd57;  #10 
a = 8'd8; b = 8'd58;  #10 
a = 8'd8; b = 8'd59;  #10 
a = 8'd8; b = 8'd60;  #10 
a = 8'd8; b = 8'd61;  #10 
a = 8'd8; b = 8'd62;  #10 
a = 8'd8; b = 8'd63;  #10 
a = 8'd8; b = 8'd64;  #10 
a = 8'd8; b = 8'd65;  #10 
a = 8'd8; b = 8'd66;  #10 
a = 8'd8; b = 8'd67;  #10 
a = 8'd8; b = 8'd68;  #10 
a = 8'd8; b = 8'd69;  #10 
a = 8'd8; b = 8'd70;  #10 
a = 8'd8; b = 8'd71;  #10 
a = 8'd8; b = 8'd72;  #10 
a = 8'd8; b = 8'd73;  #10 
a = 8'd8; b = 8'd74;  #10 
a = 8'd8; b = 8'd75;  #10 
a = 8'd8; b = 8'd76;  #10 
a = 8'd8; b = 8'd77;  #10 
a = 8'd8; b = 8'd78;  #10 
a = 8'd8; b = 8'd79;  #10 
a = 8'd8; b = 8'd80;  #10 
a = 8'd8; b = 8'd81;  #10 
a = 8'd8; b = 8'd82;  #10 
a = 8'd8; b = 8'd83;  #10 
a = 8'd8; b = 8'd84;  #10 
a = 8'd8; b = 8'd85;  #10 
a = 8'd8; b = 8'd86;  #10 
a = 8'd8; b = 8'd87;  #10 
a = 8'd8; b = 8'd88;  #10 
a = 8'd8; b = 8'd89;  #10 
a = 8'd8; b = 8'd90;  #10 
a = 8'd8; b = 8'd91;  #10 
a = 8'd8; b = 8'd92;  #10 
a = 8'd8; b = 8'd93;  #10 
a = 8'd8; b = 8'd94;  #10 
a = 8'd8; b = 8'd95;  #10 
a = 8'd8; b = 8'd96;  #10 
a = 8'd8; b = 8'd97;  #10 
a = 8'd8; b = 8'd98;  #10 
a = 8'd8; b = 8'd99;  #10 
a = 8'd8; b = 8'd100;  #10 
a = 8'd8; b = 8'd101;  #10 
a = 8'd8; b = 8'd102;  #10 
a = 8'd8; b = 8'd103;  #10 
a = 8'd8; b = 8'd104;  #10 
a = 8'd8; b = 8'd105;  #10 
a = 8'd8; b = 8'd106;  #10 
a = 8'd8; b = 8'd107;  #10 
a = 8'd8; b = 8'd108;  #10 
a = 8'd8; b = 8'd109;  #10 
a = 8'd8; b = 8'd110;  #10 
a = 8'd8; b = 8'd111;  #10 
a = 8'd8; b = 8'd112;  #10 
a = 8'd8; b = 8'd113;  #10 
a = 8'd8; b = 8'd114;  #10 
a = 8'd8; b = 8'd115;  #10 
a = 8'd8; b = 8'd116;  #10 
a = 8'd8; b = 8'd117;  #10 
a = 8'd8; b = 8'd118;  #10 
a = 8'd8; b = 8'd119;  #10 
a = 8'd8; b = 8'd120;  #10 
a = 8'd8; b = 8'd121;  #10 
a = 8'd8; b = 8'd122;  #10 
a = 8'd8; b = 8'd123;  #10 
a = 8'd8; b = 8'd124;  #10 
a = 8'd8; b = 8'd125;  #10 
a = 8'd8; b = 8'd126;  #10 
a = 8'd8; b = 8'd127;  #10 
a = 8'd8; b = 8'd128;  #10 
a = 8'd8; b = 8'd129;  #10 
a = 8'd8; b = 8'd130;  #10 
a = 8'd8; b = 8'd131;  #10 
a = 8'd8; b = 8'd132;  #10 
a = 8'd8; b = 8'd133;  #10 
a = 8'd8; b = 8'd134;  #10 
a = 8'd8; b = 8'd135;  #10 
a = 8'd8; b = 8'd136;  #10 
a = 8'd8; b = 8'd137;  #10 
a = 8'd8; b = 8'd138;  #10 
a = 8'd8; b = 8'd139;  #10 
a = 8'd8; b = 8'd140;  #10 
a = 8'd8; b = 8'd141;  #10 
a = 8'd8; b = 8'd142;  #10 
a = 8'd8; b = 8'd143;  #10 
a = 8'd8; b = 8'd144;  #10 
a = 8'd8; b = 8'd145;  #10 
a = 8'd8; b = 8'd146;  #10 
a = 8'd8; b = 8'd147;  #10 
a = 8'd8; b = 8'd148;  #10 
a = 8'd8; b = 8'd149;  #10 
a = 8'd8; b = 8'd150;  #10 
a = 8'd8; b = 8'd151;  #10 
a = 8'd8; b = 8'd152;  #10 
a = 8'd8; b = 8'd153;  #10 
a = 8'd8; b = 8'd154;  #10 
a = 8'd8; b = 8'd155;  #10 
a = 8'd8; b = 8'd156;  #10 
a = 8'd8; b = 8'd157;  #10 
a = 8'd8; b = 8'd158;  #10 
a = 8'd8; b = 8'd159;  #10 
a = 8'd8; b = 8'd160;  #10 
a = 8'd8; b = 8'd161;  #10 
a = 8'd8; b = 8'd162;  #10 
a = 8'd8; b = 8'd163;  #10 
a = 8'd8; b = 8'd164;  #10 
a = 8'd8; b = 8'd165;  #10 
a = 8'd8; b = 8'd166;  #10 
a = 8'd8; b = 8'd167;  #10 
a = 8'd8; b = 8'd168;  #10 
a = 8'd8; b = 8'd169;  #10 
a = 8'd8; b = 8'd170;  #10 
a = 8'd8; b = 8'd171;  #10 
a = 8'd8; b = 8'd172;  #10 
a = 8'd8; b = 8'd173;  #10 
a = 8'd8; b = 8'd174;  #10 
a = 8'd8; b = 8'd175;  #10 
a = 8'd8; b = 8'd176;  #10 
a = 8'd8; b = 8'd177;  #10 
a = 8'd8; b = 8'd178;  #10 
a = 8'd8; b = 8'd179;  #10 
a = 8'd8; b = 8'd180;  #10 
a = 8'd8; b = 8'd181;  #10 
a = 8'd8; b = 8'd182;  #10 
a = 8'd8; b = 8'd183;  #10 
a = 8'd8; b = 8'd184;  #10 
a = 8'd8; b = 8'd185;  #10 
a = 8'd8; b = 8'd186;  #10 
a = 8'd8; b = 8'd187;  #10 
a = 8'd8; b = 8'd188;  #10 
a = 8'd8; b = 8'd189;  #10 
a = 8'd8; b = 8'd190;  #10 
a = 8'd8; b = 8'd191;  #10 
a = 8'd8; b = 8'd192;  #10 
a = 8'd8; b = 8'd193;  #10 
a = 8'd8; b = 8'd194;  #10 
a = 8'd8; b = 8'd195;  #10 
a = 8'd8; b = 8'd196;  #10 
a = 8'd8; b = 8'd197;  #10 
a = 8'd8; b = 8'd198;  #10 
a = 8'd8; b = 8'd199;  #10 
a = 8'd8; b = 8'd200;  #10 
a = 8'd8; b = 8'd201;  #10 
a = 8'd8; b = 8'd202;  #10 
a = 8'd8; b = 8'd203;  #10 
a = 8'd8; b = 8'd204;  #10 
a = 8'd8; b = 8'd205;  #10 
a = 8'd8; b = 8'd206;  #10 
a = 8'd8; b = 8'd207;  #10 
a = 8'd8; b = 8'd208;  #10 
a = 8'd8; b = 8'd209;  #10 
a = 8'd8; b = 8'd210;  #10 
a = 8'd8; b = 8'd211;  #10 
a = 8'd8; b = 8'd212;  #10 
a = 8'd8; b = 8'd213;  #10 
a = 8'd8; b = 8'd214;  #10 
a = 8'd8; b = 8'd215;  #10 
a = 8'd8; b = 8'd216;  #10 
a = 8'd8; b = 8'd217;  #10 
a = 8'd8; b = 8'd218;  #10 
a = 8'd8; b = 8'd219;  #10 
a = 8'd8; b = 8'd220;  #10 
a = 8'd8; b = 8'd221;  #10 
a = 8'd8; b = 8'd222;  #10 
a = 8'd8; b = 8'd223;  #10 
a = 8'd8; b = 8'd224;  #10 
a = 8'd8; b = 8'd225;  #10 
a = 8'd8; b = 8'd226;  #10 
a = 8'd8; b = 8'd227;  #10 
a = 8'd8; b = 8'd228;  #10 
a = 8'd8; b = 8'd229;  #10 
a = 8'd8; b = 8'd230;  #10 
a = 8'd8; b = 8'd231;  #10 
a = 8'd8; b = 8'd232;  #10 
a = 8'd8; b = 8'd233;  #10 
a = 8'd8; b = 8'd234;  #10 
a = 8'd8; b = 8'd235;  #10 
a = 8'd8; b = 8'd236;  #10 
a = 8'd8; b = 8'd237;  #10 
a = 8'd8; b = 8'd238;  #10 
a = 8'd8; b = 8'd239;  #10 
a = 8'd8; b = 8'd240;  #10 
a = 8'd8; b = 8'd241;  #10 
a = 8'd8; b = 8'd242;  #10 
a = 8'd8; b = 8'd243;  #10 
a = 8'd8; b = 8'd244;  #10 
a = 8'd8; b = 8'd245;  #10 
a = 8'd8; b = 8'd246;  #10 
a = 8'd8; b = 8'd247;  #10 
a = 8'd8; b = 8'd248;  #10 
a = 8'd8; b = 8'd249;  #10 
a = 8'd8; b = 8'd250;  #10 
a = 8'd8; b = 8'd251;  #10 
a = 8'd8; b = 8'd252;  #10 
a = 8'd8; b = 8'd253;  #10 
a = 8'd8; b = 8'd254;  #10 
a = 8'd8; b = 8'd255;  #10 
a = 8'd9; b = 8'd0;  #10 
a = 8'd9; b = 8'd1;  #10 
a = 8'd9; b = 8'd2;  #10 
a = 8'd9; b = 8'd3;  #10 
a = 8'd9; b = 8'd4;  #10 
a = 8'd9; b = 8'd5;  #10 
a = 8'd9; b = 8'd6;  #10 
a = 8'd9; b = 8'd7;  #10 
a = 8'd9; b = 8'd8;  #10 
a = 8'd9; b = 8'd9;  #10 
a = 8'd9; b = 8'd10;  #10 
a = 8'd9; b = 8'd11;  #10 
a = 8'd9; b = 8'd12;  #10 
a = 8'd9; b = 8'd13;  #10 
a = 8'd9; b = 8'd14;  #10 
a = 8'd9; b = 8'd15;  #10 
a = 8'd9; b = 8'd16;  #10 
a = 8'd9; b = 8'd17;  #10 
a = 8'd9; b = 8'd18;  #10 
a = 8'd9; b = 8'd19;  #10 
a = 8'd9; b = 8'd20;  #10 
a = 8'd9; b = 8'd21;  #10 
a = 8'd9; b = 8'd22;  #10 
a = 8'd9; b = 8'd23;  #10 
a = 8'd9; b = 8'd24;  #10 
a = 8'd9; b = 8'd25;  #10 
a = 8'd9; b = 8'd26;  #10 
a = 8'd9; b = 8'd27;  #10 
a = 8'd9; b = 8'd28;  #10 
a = 8'd9; b = 8'd29;  #10 
a = 8'd9; b = 8'd30;  #10 
a = 8'd9; b = 8'd31;  #10 
a = 8'd9; b = 8'd32;  #10 
a = 8'd9; b = 8'd33;  #10 
a = 8'd9; b = 8'd34;  #10 
a = 8'd9; b = 8'd35;  #10 
a = 8'd9; b = 8'd36;  #10 
a = 8'd9; b = 8'd37;  #10 
a = 8'd9; b = 8'd38;  #10 
a = 8'd9; b = 8'd39;  #10 
a = 8'd9; b = 8'd40;  #10 
a = 8'd9; b = 8'd41;  #10 
a = 8'd9; b = 8'd42;  #10 
a = 8'd9; b = 8'd43;  #10 
a = 8'd9; b = 8'd44;  #10 
a = 8'd9; b = 8'd45;  #10 
a = 8'd9; b = 8'd46;  #10 
a = 8'd9; b = 8'd47;  #10 
a = 8'd9; b = 8'd48;  #10 
a = 8'd9; b = 8'd49;  #10 
a = 8'd9; b = 8'd50;  #10 
a = 8'd9; b = 8'd51;  #10 
a = 8'd9; b = 8'd52;  #10 
a = 8'd9; b = 8'd53;  #10 
a = 8'd9; b = 8'd54;  #10 
a = 8'd9; b = 8'd55;  #10 
a = 8'd9; b = 8'd56;  #10 
a = 8'd9; b = 8'd57;  #10 
a = 8'd9; b = 8'd58;  #10 
a = 8'd9; b = 8'd59;  #10 
a = 8'd9; b = 8'd60;  #10 
a = 8'd9; b = 8'd61;  #10 
a = 8'd9; b = 8'd62;  #10 
a = 8'd9; b = 8'd63;  #10 
a = 8'd9; b = 8'd64;  #10 
a = 8'd9; b = 8'd65;  #10 
a = 8'd9; b = 8'd66;  #10 
a = 8'd9; b = 8'd67;  #10 
a = 8'd9; b = 8'd68;  #10 
a = 8'd9; b = 8'd69;  #10 
a = 8'd9; b = 8'd70;  #10 
a = 8'd9; b = 8'd71;  #10 
a = 8'd9; b = 8'd72;  #10 
a = 8'd9; b = 8'd73;  #10 
a = 8'd9; b = 8'd74;  #10 
a = 8'd9; b = 8'd75;  #10 
a = 8'd9; b = 8'd76;  #10 
a = 8'd9; b = 8'd77;  #10 
a = 8'd9; b = 8'd78;  #10 
a = 8'd9; b = 8'd79;  #10 
a = 8'd9; b = 8'd80;  #10 
a = 8'd9; b = 8'd81;  #10 
a = 8'd9; b = 8'd82;  #10 
a = 8'd9; b = 8'd83;  #10 
a = 8'd9; b = 8'd84;  #10 
a = 8'd9; b = 8'd85;  #10 
a = 8'd9; b = 8'd86;  #10 
a = 8'd9; b = 8'd87;  #10 
a = 8'd9; b = 8'd88;  #10 
a = 8'd9; b = 8'd89;  #10 
a = 8'd9; b = 8'd90;  #10 
a = 8'd9; b = 8'd91;  #10 
a = 8'd9; b = 8'd92;  #10 
a = 8'd9; b = 8'd93;  #10 
a = 8'd9; b = 8'd94;  #10 
a = 8'd9; b = 8'd95;  #10 
a = 8'd9; b = 8'd96;  #10 
a = 8'd9; b = 8'd97;  #10 
a = 8'd9; b = 8'd98;  #10 
a = 8'd9; b = 8'd99;  #10 
a = 8'd9; b = 8'd100;  #10 
a = 8'd9; b = 8'd101;  #10 
a = 8'd9; b = 8'd102;  #10 
a = 8'd9; b = 8'd103;  #10 
a = 8'd9; b = 8'd104;  #10 
a = 8'd9; b = 8'd105;  #10 
a = 8'd9; b = 8'd106;  #10 
a = 8'd9; b = 8'd107;  #10 
a = 8'd9; b = 8'd108;  #10 
a = 8'd9; b = 8'd109;  #10 
a = 8'd9; b = 8'd110;  #10 
a = 8'd9; b = 8'd111;  #10 
a = 8'd9; b = 8'd112;  #10 
a = 8'd9; b = 8'd113;  #10 
a = 8'd9; b = 8'd114;  #10 
a = 8'd9; b = 8'd115;  #10 
a = 8'd9; b = 8'd116;  #10 
a = 8'd9; b = 8'd117;  #10 
a = 8'd9; b = 8'd118;  #10 
a = 8'd9; b = 8'd119;  #10 
a = 8'd9; b = 8'd120;  #10 
a = 8'd9; b = 8'd121;  #10 
a = 8'd9; b = 8'd122;  #10 
a = 8'd9; b = 8'd123;  #10 
a = 8'd9; b = 8'd124;  #10 
a = 8'd9; b = 8'd125;  #10 
a = 8'd9; b = 8'd126;  #10 
a = 8'd9; b = 8'd127;  #10 
a = 8'd9; b = 8'd128;  #10 
a = 8'd9; b = 8'd129;  #10 
a = 8'd9; b = 8'd130;  #10 
a = 8'd9; b = 8'd131;  #10 
a = 8'd9; b = 8'd132;  #10 
a = 8'd9; b = 8'd133;  #10 
a = 8'd9; b = 8'd134;  #10 
a = 8'd9; b = 8'd135;  #10 
a = 8'd9; b = 8'd136;  #10 
a = 8'd9; b = 8'd137;  #10 
a = 8'd9; b = 8'd138;  #10 
a = 8'd9; b = 8'd139;  #10 
a = 8'd9; b = 8'd140;  #10 
a = 8'd9; b = 8'd141;  #10 
a = 8'd9; b = 8'd142;  #10 
a = 8'd9; b = 8'd143;  #10 
a = 8'd9; b = 8'd144;  #10 
a = 8'd9; b = 8'd145;  #10 
a = 8'd9; b = 8'd146;  #10 
a = 8'd9; b = 8'd147;  #10 
a = 8'd9; b = 8'd148;  #10 
a = 8'd9; b = 8'd149;  #10 
a = 8'd9; b = 8'd150;  #10 
a = 8'd9; b = 8'd151;  #10 
a = 8'd9; b = 8'd152;  #10 
a = 8'd9; b = 8'd153;  #10 
a = 8'd9; b = 8'd154;  #10 
a = 8'd9; b = 8'd155;  #10 
a = 8'd9; b = 8'd156;  #10 
a = 8'd9; b = 8'd157;  #10 
a = 8'd9; b = 8'd158;  #10 
a = 8'd9; b = 8'd159;  #10 
a = 8'd9; b = 8'd160;  #10 
a = 8'd9; b = 8'd161;  #10 
a = 8'd9; b = 8'd162;  #10 
a = 8'd9; b = 8'd163;  #10 
a = 8'd9; b = 8'd164;  #10 
a = 8'd9; b = 8'd165;  #10 
a = 8'd9; b = 8'd166;  #10 
a = 8'd9; b = 8'd167;  #10 
a = 8'd9; b = 8'd168;  #10 
a = 8'd9; b = 8'd169;  #10 
a = 8'd9; b = 8'd170;  #10 
a = 8'd9; b = 8'd171;  #10 
a = 8'd9; b = 8'd172;  #10 
a = 8'd9; b = 8'd173;  #10 
a = 8'd9; b = 8'd174;  #10 
a = 8'd9; b = 8'd175;  #10 
a = 8'd9; b = 8'd176;  #10 
a = 8'd9; b = 8'd177;  #10 
a = 8'd9; b = 8'd178;  #10 
a = 8'd9; b = 8'd179;  #10 
a = 8'd9; b = 8'd180;  #10 
a = 8'd9; b = 8'd181;  #10 
a = 8'd9; b = 8'd182;  #10 
a = 8'd9; b = 8'd183;  #10 
a = 8'd9; b = 8'd184;  #10 
a = 8'd9; b = 8'd185;  #10 
a = 8'd9; b = 8'd186;  #10 
a = 8'd9; b = 8'd187;  #10 
a = 8'd9; b = 8'd188;  #10 
a = 8'd9; b = 8'd189;  #10 
a = 8'd9; b = 8'd190;  #10 
a = 8'd9; b = 8'd191;  #10 
a = 8'd9; b = 8'd192;  #10 
a = 8'd9; b = 8'd193;  #10 
a = 8'd9; b = 8'd194;  #10 
a = 8'd9; b = 8'd195;  #10 
a = 8'd9; b = 8'd196;  #10 
a = 8'd9; b = 8'd197;  #10 
a = 8'd9; b = 8'd198;  #10 
a = 8'd9; b = 8'd199;  #10 
a = 8'd9; b = 8'd200;  #10 
a = 8'd9; b = 8'd201;  #10 
a = 8'd9; b = 8'd202;  #10 
a = 8'd9; b = 8'd203;  #10 
a = 8'd9; b = 8'd204;  #10 
a = 8'd9; b = 8'd205;  #10 
a = 8'd9; b = 8'd206;  #10 
a = 8'd9; b = 8'd207;  #10 
a = 8'd9; b = 8'd208;  #10 
a = 8'd9; b = 8'd209;  #10 
a = 8'd9; b = 8'd210;  #10 
a = 8'd9; b = 8'd211;  #10 
a = 8'd9; b = 8'd212;  #10 
a = 8'd9; b = 8'd213;  #10 
a = 8'd9; b = 8'd214;  #10 
a = 8'd9; b = 8'd215;  #10 
a = 8'd9; b = 8'd216;  #10 
a = 8'd9; b = 8'd217;  #10 
a = 8'd9; b = 8'd218;  #10 
a = 8'd9; b = 8'd219;  #10 
a = 8'd9; b = 8'd220;  #10 
a = 8'd9; b = 8'd221;  #10 
a = 8'd9; b = 8'd222;  #10 
a = 8'd9; b = 8'd223;  #10 
a = 8'd9; b = 8'd224;  #10 
a = 8'd9; b = 8'd225;  #10 
a = 8'd9; b = 8'd226;  #10 
a = 8'd9; b = 8'd227;  #10 
a = 8'd9; b = 8'd228;  #10 
a = 8'd9; b = 8'd229;  #10 
a = 8'd9; b = 8'd230;  #10 
a = 8'd9; b = 8'd231;  #10 
a = 8'd9; b = 8'd232;  #10 
a = 8'd9; b = 8'd233;  #10 
a = 8'd9; b = 8'd234;  #10 
a = 8'd9; b = 8'd235;  #10 
a = 8'd9; b = 8'd236;  #10 
a = 8'd9; b = 8'd237;  #10 
a = 8'd9; b = 8'd238;  #10 
a = 8'd9; b = 8'd239;  #10 
a = 8'd9; b = 8'd240;  #10 
a = 8'd9; b = 8'd241;  #10 
a = 8'd9; b = 8'd242;  #10 
a = 8'd9; b = 8'd243;  #10 
a = 8'd9; b = 8'd244;  #10 
a = 8'd9; b = 8'd245;  #10 
a = 8'd9; b = 8'd246;  #10 
a = 8'd9; b = 8'd247;  #10 
a = 8'd9; b = 8'd248;  #10 
a = 8'd9; b = 8'd249;  #10 
a = 8'd9; b = 8'd250;  #10 
a = 8'd9; b = 8'd251;  #10 
a = 8'd9; b = 8'd252;  #10 
a = 8'd9; b = 8'd253;  #10 
a = 8'd9; b = 8'd254;  #10 
a = 8'd9; b = 8'd255;  #10 
a = 8'd10; b = 8'd0;  #10 
a = 8'd10; b = 8'd1;  #10 
a = 8'd10; b = 8'd2;  #10 
a = 8'd10; b = 8'd3;  #10 
a = 8'd10; b = 8'd4;  #10 
a = 8'd10; b = 8'd5;  #10 
a = 8'd10; b = 8'd6;  #10 
a = 8'd10; b = 8'd7;  #10 
a = 8'd10; b = 8'd8;  #10 
a = 8'd10; b = 8'd9;  #10 
a = 8'd10; b = 8'd10;  #10 
a = 8'd10; b = 8'd11;  #10 
a = 8'd10; b = 8'd12;  #10 
a = 8'd10; b = 8'd13;  #10 
a = 8'd10; b = 8'd14;  #10 
a = 8'd10; b = 8'd15;  #10 
a = 8'd10; b = 8'd16;  #10 
a = 8'd10; b = 8'd17;  #10 
a = 8'd10; b = 8'd18;  #10 
a = 8'd10; b = 8'd19;  #10 
a = 8'd10; b = 8'd20;  #10 
a = 8'd10; b = 8'd21;  #10 
a = 8'd10; b = 8'd22;  #10 
a = 8'd10; b = 8'd23;  #10 
a = 8'd10; b = 8'd24;  #10 
a = 8'd10; b = 8'd25;  #10 
a = 8'd10; b = 8'd26;  #10 
a = 8'd10; b = 8'd27;  #10 
a = 8'd10; b = 8'd28;  #10 
a = 8'd10; b = 8'd29;  #10 
a = 8'd10; b = 8'd30;  #10 
a = 8'd10; b = 8'd31;  #10 
a = 8'd10; b = 8'd32;  #10 
a = 8'd10; b = 8'd33;  #10 
a = 8'd10; b = 8'd34;  #10 
a = 8'd10; b = 8'd35;  #10 
a = 8'd10; b = 8'd36;  #10 
a = 8'd10; b = 8'd37;  #10 
a = 8'd10; b = 8'd38;  #10 
a = 8'd10; b = 8'd39;  #10 
a = 8'd10; b = 8'd40;  #10 
a = 8'd10; b = 8'd41;  #10 
a = 8'd10; b = 8'd42;  #10 
a = 8'd10; b = 8'd43;  #10 
a = 8'd10; b = 8'd44;  #10 
a = 8'd10; b = 8'd45;  #10 
a = 8'd10; b = 8'd46;  #10 
a = 8'd10; b = 8'd47;  #10 
a = 8'd10; b = 8'd48;  #10 
a = 8'd10; b = 8'd49;  #10 
a = 8'd10; b = 8'd50;  #10 
a = 8'd10; b = 8'd51;  #10 
a = 8'd10; b = 8'd52;  #10 
a = 8'd10; b = 8'd53;  #10 
a = 8'd10; b = 8'd54;  #10 
a = 8'd10; b = 8'd55;  #10 
a = 8'd10; b = 8'd56;  #10 
a = 8'd10; b = 8'd57;  #10 
a = 8'd10; b = 8'd58;  #10 
a = 8'd10; b = 8'd59;  #10 
a = 8'd10; b = 8'd60;  #10 
a = 8'd10; b = 8'd61;  #10 
a = 8'd10; b = 8'd62;  #10 
a = 8'd10; b = 8'd63;  #10 
a = 8'd10; b = 8'd64;  #10 
a = 8'd10; b = 8'd65;  #10 
a = 8'd10; b = 8'd66;  #10 
a = 8'd10; b = 8'd67;  #10 
a = 8'd10; b = 8'd68;  #10 
a = 8'd10; b = 8'd69;  #10 
a = 8'd10; b = 8'd70;  #10 
a = 8'd10; b = 8'd71;  #10 
a = 8'd10; b = 8'd72;  #10 
a = 8'd10; b = 8'd73;  #10 
a = 8'd10; b = 8'd74;  #10 
a = 8'd10; b = 8'd75;  #10 
a = 8'd10; b = 8'd76;  #10 
a = 8'd10; b = 8'd77;  #10 
a = 8'd10; b = 8'd78;  #10 
a = 8'd10; b = 8'd79;  #10 
a = 8'd10; b = 8'd80;  #10 
a = 8'd10; b = 8'd81;  #10 
a = 8'd10; b = 8'd82;  #10 
a = 8'd10; b = 8'd83;  #10 
a = 8'd10; b = 8'd84;  #10 
a = 8'd10; b = 8'd85;  #10 
a = 8'd10; b = 8'd86;  #10 
a = 8'd10; b = 8'd87;  #10 
a = 8'd10; b = 8'd88;  #10 
a = 8'd10; b = 8'd89;  #10 
a = 8'd10; b = 8'd90;  #10 
a = 8'd10; b = 8'd91;  #10 
a = 8'd10; b = 8'd92;  #10 
a = 8'd10; b = 8'd93;  #10 
a = 8'd10; b = 8'd94;  #10 
a = 8'd10; b = 8'd95;  #10 
a = 8'd10; b = 8'd96;  #10 
a = 8'd10; b = 8'd97;  #10 
a = 8'd10; b = 8'd98;  #10 
a = 8'd10; b = 8'd99;  #10 
a = 8'd10; b = 8'd100;  #10 
a = 8'd10; b = 8'd101;  #10 
a = 8'd10; b = 8'd102;  #10 
a = 8'd10; b = 8'd103;  #10 
a = 8'd10; b = 8'd104;  #10 
a = 8'd10; b = 8'd105;  #10 
a = 8'd10; b = 8'd106;  #10 
a = 8'd10; b = 8'd107;  #10 
a = 8'd10; b = 8'd108;  #10 
a = 8'd10; b = 8'd109;  #10 
a = 8'd10; b = 8'd110;  #10 
a = 8'd10; b = 8'd111;  #10 
a = 8'd10; b = 8'd112;  #10 
a = 8'd10; b = 8'd113;  #10 
a = 8'd10; b = 8'd114;  #10 
a = 8'd10; b = 8'd115;  #10 
a = 8'd10; b = 8'd116;  #10 
a = 8'd10; b = 8'd117;  #10 
a = 8'd10; b = 8'd118;  #10 
a = 8'd10; b = 8'd119;  #10 
a = 8'd10; b = 8'd120;  #10 
a = 8'd10; b = 8'd121;  #10 
a = 8'd10; b = 8'd122;  #10 
a = 8'd10; b = 8'd123;  #10 
a = 8'd10; b = 8'd124;  #10 
a = 8'd10; b = 8'd125;  #10 
a = 8'd10; b = 8'd126;  #10 
a = 8'd10; b = 8'd127;  #10 
a = 8'd10; b = 8'd128;  #10 
a = 8'd10; b = 8'd129;  #10 
a = 8'd10; b = 8'd130;  #10 
a = 8'd10; b = 8'd131;  #10 
a = 8'd10; b = 8'd132;  #10 
a = 8'd10; b = 8'd133;  #10 
a = 8'd10; b = 8'd134;  #10 
a = 8'd10; b = 8'd135;  #10 
a = 8'd10; b = 8'd136;  #10 
a = 8'd10; b = 8'd137;  #10 
a = 8'd10; b = 8'd138;  #10 
a = 8'd10; b = 8'd139;  #10 
a = 8'd10; b = 8'd140;  #10 
a = 8'd10; b = 8'd141;  #10 
a = 8'd10; b = 8'd142;  #10 
a = 8'd10; b = 8'd143;  #10 
a = 8'd10; b = 8'd144;  #10 
a = 8'd10; b = 8'd145;  #10 
a = 8'd10; b = 8'd146;  #10 
a = 8'd10; b = 8'd147;  #10 
a = 8'd10; b = 8'd148;  #10 
a = 8'd10; b = 8'd149;  #10 
a = 8'd10; b = 8'd150;  #10 
a = 8'd10; b = 8'd151;  #10 
a = 8'd10; b = 8'd152;  #10 
a = 8'd10; b = 8'd153;  #10 
a = 8'd10; b = 8'd154;  #10 
a = 8'd10; b = 8'd155;  #10 
a = 8'd10; b = 8'd156;  #10 
a = 8'd10; b = 8'd157;  #10 
a = 8'd10; b = 8'd158;  #10 
a = 8'd10; b = 8'd159;  #10 
a = 8'd10; b = 8'd160;  #10 
a = 8'd10; b = 8'd161;  #10 
a = 8'd10; b = 8'd162;  #10 
a = 8'd10; b = 8'd163;  #10 
a = 8'd10; b = 8'd164;  #10 
a = 8'd10; b = 8'd165;  #10 
a = 8'd10; b = 8'd166;  #10 
a = 8'd10; b = 8'd167;  #10 
a = 8'd10; b = 8'd168;  #10 
a = 8'd10; b = 8'd169;  #10 
a = 8'd10; b = 8'd170;  #10 
a = 8'd10; b = 8'd171;  #10 
a = 8'd10; b = 8'd172;  #10 
a = 8'd10; b = 8'd173;  #10 
a = 8'd10; b = 8'd174;  #10 
a = 8'd10; b = 8'd175;  #10 
a = 8'd10; b = 8'd176;  #10 
a = 8'd10; b = 8'd177;  #10 
a = 8'd10; b = 8'd178;  #10 
a = 8'd10; b = 8'd179;  #10 
a = 8'd10; b = 8'd180;  #10 
a = 8'd10; b = 8'd181;  #10 
a = 8'd10; b = 8'd182;  #10 
a = 8'd10; b = 8'd183;  #10 
a = 8'd10; b = 8'd184;  #10 
a = 8'd10; b = 8'd185;  #10 
a = 8'd10; b = 8'd186;  #10 
a = 8'd10; b = 8'd187;  #10 
a = 8'd10; b = 8'd188;  #10 
a = 8'd10; b = 8'd189;  #10 
a = 8'd10; b = 8'd190;  #10 
a = 8'd10; b = 8'd191;  #10 
a = 8'd10; b = 8'd192;  #10 
a = 8'd10; b = 8'd193;  #10 
a = 8'd10; b = 8'd194;  #10 
a = 8'd10; b = 8'd195;  #10 
a = 8'd10; b = 8'd196;  #10 
a = 8'd10; b = 8'd197;  #10 
a = 8'd10; b = 8'd198;  #10 
a = 8'd10; b = 8'd199;  #10 
a = 8'd10; b = 8'd200;  #10 
a = 8'd10; b = 8'd201;  #10 
a = 8'd10; b = 8'd202;  #10 
a = 8'd10; b = 8'd203;  #10 
a = 8'd10; b = 8'd204;  #10 
a = 8'd10; b = 8'd205;  #10 
a = 8'd10; b = 8'd206;  #10 
a = 8'd10; b = 8'd207;  #10 
a = 8'd10; b = 8'd208;  #10 
a = 8'd10; b = 8'd209;  #10 
a = 8'd10; b = 8'd210;  #10 
a = 8'd10; b = 8'd211;  #10 
a = 8'd10; b = 8'd212;  #10 
a = 8'd10; b = 8'd213;  #10 
a = 8'd10; b = 8'd214;  #10 
a = 8'd10; b = 8'd215;  #10 
a = 8'd10; b = 8'd216;  #10 
a = 8'd10; b = 8'd217;  #10 
a = 8'd10; b = 8'd218;  #10 
a = 8'd10; b = 8'd219;  #10 
a = 8'd10; b = 8'd220;  #10 
a = 8'd10; b = 8'd221;  #10 
a = 8'd10; b = 8'd222;  #10 
a = 8'd10; b = 8'd223;  #10 
a = 8'd10; b = 8'd224;  #10 
a = 8'd10; b = 8'd225;  #10 
a = 8'd10; b = 8'd226;  #10 
a = 8'd10; b = 8'd227;  #10 
a = 8'd10; b = 8'd228;  #10 
a = 8'd10; b = 8'd229;  #10 
a = 8'd10; b = 8'd230;  #10 
a = 8'd10; b = 8'd231;  #10 
a = 8'd10; b = 8'd232;  #10 
a = 8'd10; b = 8'd233;  #10 
a = 8'd10; b = 8'd234;  #10 
a = 8'd10; b = 8'd235;  #10 
a = 8'd10; b = 8'd236;  #10 
a = 8'd10; b = 8'd237;  #10 
a = 8'd10; b = 8'd238;  #10 
a = 8'd10; b = 8'd239;  #10 
a = 8'd10; b = 8'd240;  #10 
a = 8'd10; b = 8'd241;  #10 
a = 8'd10; b = 8'd242;  #10 
a = 8'd10; b = 8'd243;  #10 
a = 8'd10; b = 8'd244;  #10 
a = 8'd10; b = 8'd245;  #10 
a = 8'd10; b = 8'd246;  #10 
a = 8'd10; b = 8'd247;  #10 
a = 8'd10; b = 8'd248;  #10 
a = 8'd10; b = 8'd249;  #10 
a = 8'd10; b = 8'd250;  #10 
a = 8'd10; b = 8'd251;  #10 
a = 8'd10; b = 8'd252;  #10 
a = 8'd10; b = 8'd253;  #10 
a = 8'd10; b = 8'd254;  #10 
a = 8'd10; b = 8'd255;  #10 
a = 8'd11; b = 8'd0;  #10 
a = 8'd11; b = 8'd1;  #10 
a = 8'd11; b = 8'd2;  #10 
a = 8'd11; b = 8'd3;  #10 
a = 8'd11; b = 8'd4;  #10 
a = 8'd11; b = 8'd5;  #10 
a = 8'd11; b = 8'd6;  #10 
a = 8'd11; b = 8'd7;  #10 
a = 8'd11; b = 8'd8;  #10 
a = 8'd11; b = 8'd9;  #10 
a = 8'd11; b = 8'd10;  #10 
a = 8'd11; b = 8'd11;  #10 
a = 8'd11; b = 8'd12;  #10 
a = 8'd11; b = 8'd13;  #10 
a = 8'd11; b = 8'd14;  #10 
a = 8'd11; b = 8'd15;  #10 
a = 8'd11; b = 8'd16;  #10 
a = 8'd11; b = 8'd17;  #10 
a = 8'd11; b = 8'd18;  #10 
a = 8'd11; b = 8'd19;  #10 
a = 8'd11; b = 8'd20;  #10 
a = 8'd11; b = 8'd21;  #10 
a = 8'd11; b = 8'd22;  #10 
a = 8'd11; b = 8'd23;  #10 
a = 8'd11; b = 8'd24;  #10 
a = 8'd11; b = 8'd25;  #10 
a = 8'd11; b = 8'd26;  #10 
a = 8'd11; b = 8'd27;  #10 
a = 8'd11; b = 8'd28;  #10 
a = 8'd11; b = 8'd29;  #10 
a = 8'd11; b = 8'd30;  #10 
a = 8'd11; b = 8'd31;  #10 
a = 8'd11; b = 8'd32;  #10 
a = 8'd11; b = 8'd33;  #10 
a = 8'd11; b = 8'd34;  #10 
a = 8'd11; b = 8'd35;  #10 
a = 8'd11; b = 8'd36;  #10 
a = 8'd11; b = 8'd37;  #10 
a = 8'd11; b = 8'd38;  #10 
a = 8'd11; b = 8'd39;  #10 
a = 8'd11; b = 8'd40;  #10 
a = 8'd11; b = 8'd41;  #10 
a = 8'd11; b = 8'd42;  #10 
a = 8'd11; b = 8'd43;  #10 
a = 8'd11; b = 8'd44;  #10 
a = 8'd11; b = 8'd45;  #10 
a = 8'd11; b = 8'd46;  #10 
a = 8'd11; b = 8'd47;  #10 
a = 8'd11; b = 8'd48;  #10 
a = 8'd11; b = 8'd49;  #10 
a = 8'd11; b = 8'd50;  #10 
a = 8'd11; b = 8'd51;  #10 
a = 8'd11; b = 8'd52;  #10 
a = 8'd11; b = 8'd53;  #10 
a = 8'd11; b = 8'd54;  #10 
a = 8'd11; b = 8'd55;  #10 
a = 8'd11; b = 8'd56;  #10 
a = 8'd11; b = 8'd57;  #10 
a = 8'd11; b = 8'd58;  #10 
a = 8'd11; b = 8'd59;  #10 
a = 8'd11; b = 8'd60;  #10 
a = 8'd11; b = 8'd61;  #10 
a = 8'd11; b = 8'd62;  #10 
a = 8'd11; b = 8'd63;  #10 
a = 8'd11; b = 8'd64;  #10 
a = 8'd11; b = 8'd65;  #10 
a = 8'd11; b = 8'd66;  #10 
a = 8'd11; b = 8'd67;  #10 
a = 8'd11; b = 8'd68;  #10 
a = 8'd11; b = 8'd69;  #10 
a = 8'd11; b = 8'd70;  #10 
a = 8'd11; b = 8'd71;  #10 
a = 8'd11; b = 8'd72;  #10 
a = 8'd11; b = 8'd73;  #10 
a = 8'd11; b = 8'd74;  #10 
a = 8'd11; b = 8'd75;  #10 
a = 8'd11; b = 8'd76;  #10 
a = 8'd11; b = 8'd77;  #10 
a = 8'd11; b = 8'd78;  #10 
a = 8'd11; b = 8'd79;  #10 
a = 8'd11; b = 8'd80;  #10 
a = 8'd11; b = 8'd81;  #10 
a = 8'd11; b = 8'd82;  #10 
a = 8'd11; b = 8'd83;  #10 
a = 8'd11; b = 8'd84;  #10 
a = 8'd11; b = 8'd85;  #10 
a = 8'd11; b = 8'd86;  #10 
a = 8'd11; b = 8'd87;  #10 
a = 8'd11; b = 8'd88;  #10 
a = 8'd11; b = 8'd89;  #10 
a = 8'd11; b = 8'd90;  #10 
a = 8'd11; b = 8'd91;  #10 
a = 8'd11; b = 8'd92;  #10 
a = 8'd11; b = 8'd93;  #10 
a = 8'd11; b = 8'd94;  #10 
a = 8'd11; b = 8'd95;  #10 
a = 8'd11; b = 8'd96;  #10 
a = 8'd11; b = 8'd97;  #10 
a = 8'd11; b = 8'd98;  #10 
a = 8'd11; b = 8'd99;  #10 
a = 8'd11; b = 8'd100;  #10 
a = 8'd11; b = 8'd101;  #10 
a = 8'd11; b = 8'd102;  #10 
a = 8'd11; b = 8'd103;  #10 
a = 8'd11; b = 8'd104;  #10 
a = 8'd11; b = 8'd105;  #10 
a = 8'd11; b = 8'd106;  #10 
a = 8'd11; b = 8'd107;  #10 
a = 8'd11; b = 8'd108;  #10 
a = 8'd11; b = 8'd109;  #10 
a = 8'd11; b = 8'd110;  #10 
a = 8'd11; b = 8'd111;  #10 
a = 8'd11; b = 8'd112;  #10 
a = 8'd11; b = 8'd113;  #10 
a = 8'd11; b = 8'd114;  #10 
a = 8'd11; b = 8'd115;  #10 
a = 8'd11; b = 8'd116;  #10 
a = 8'd11; b = 8'd117;  #10 
a = 8'd11; b = 8'd118;  #10 
a = 8'd11; b = 8'd119;  #10 
a = 8'd11; b = 8'd120;  #10 
a = 8'd11; b = 8'd121;  #10 
a = 8'd11; b = 8'd122;  #10 
a = 8'd11; b = 8'd123;  #10 
a = 8'd11; b = 8'd124;  #10 
a = 8'd11; b = 8'd125;  #10 
a = 8'd11; b = 8'd126;  #10 
a = 8'd11; b = 8'd127;  #10 
a = 8'd11; b = 8'd128;  #10 
a = 8'd11; b = 8'd129;  #10 
a = 8'd11; b = 8'd130;  #10 
a = 8'd11; b = 8'd131;  #10 
a = 8'd11; b = 8'd132;  #10 
a = 8'd11; b = 8'd133;  #10 
a = 8'd11; b = 8'd134;  #10 
a = 8'd11; b = 8'd135;  #10 
a = 8'd11; b = 8'd136;  #10 
a = 8'd11; b = 8'd137;  #10 
a = 8'd11; b = 8'd138;  #10 
a = 8'd11; b = 8'd139;  #10 
a = 8'd11; b = 8'd140;  #10 
a = 8'd11; b = 8'd141;  #10 
a = 8'd11; b = 8'd142;  #10 
a = 8'd11; b = 8'd143;  #10 
a = 8'd11; b = 8'd144;  #10 
a = 8'd11; b = 8'd145;  #10 
a = 8'd11; b = 8'd146;  #10 
a = 8'd11; b = 8'd147;  #10 
a = 8'd11; b = 8'd148;  #10 
a = 8'd11; b = 8'd149;  #10 
a = 8'd11; b = 8'd150;  #10 
a = 8'd11; b = 8'd151;  #10 
a = 8'd11; b = 8'd152;  #10 
a = 8'd11; b = 8'd153;  #10 
a = 8'd11; b = 8'd154;  #10 
a = 8'd11; b = 8'd155;  #10 
a = 8'd11; b = 8'd156;  #10 
a = 8'd11; b = 8'd157;  #10 
a = 8'd11; b = 8'd158;  #10 
a = 8'd11; b = 8'd159;  #10 
a = 8'd11; b = 8'd160;  #10 
a = 8'd11; b = 8'd161;  #10 
a = 8'd11; b = 8'd162;  #10 
a = 8'd11; b = 8'd163;  #10 
a = 8'd11; b = 8'd164;  #10 
a = 8'd11; b = 8'd165;  #10 
a = 8'd11; b = 8'd166;  #10 
a = 8'd11; b = 8'd167;  #10 
a = 8'd11; b = 8'd168;  #10 
a = 8'd11; b = 8'd169;  #10 
a = 8'd11; b = 8'd170;  #10 
a = 8'd11; b = 8'd171;  #10 
a = 8'd11; b = 8'd172;  #10 
a = 8'd11; b = 8'd173;  #10 
a = 8'd11; b = 8'd174;  #10 
a = 8'd11; b = 8'd175;  #10 
a = 8'd11; b = 8'd176;  #10 
a = 8'd11; b = 8'd177;  #10 
a = 8'd11; b = 8'd178;  #10 
a = 8'd11; b = 8'd179;  #10 
a = 8'd11; b = 8'd180;  #10 
a = 8'd11; b = 8'd181;  #10 
a = 8'd11; b = 8'd182;  #10 
a = 8'd11; b = 8'd183;  #10 
a = 8'd11; b = 8'd184;  #10 
a = 8'd11; b = 8'd185;  #10 
a = 8'd11; b = 8'd186;  #10 
a = 8'd11; b = 8'd187;  #10 
a = 8'd11; b = 8'd188;  #10 
a = 8'd11; b = 8'd189;  #10 
a = 8'd11; b = 8'd190;  #10 
a = 8'd11; b = 8'd191;  #10 
a = 8'd11; b = 8'd192;  #10 
a = 8'd11; b = 8'd193;  #10 
a = 8'd11; b = 8'd194;  #10 
a = 8'd11; b = 8'd195;  #10 
a = 8'd11; b = 8'd196;  #10 
a = 8'd11; b = 8'd197;  #10 
a = 8'd11; b = 8'd198;  #10 
a = 8'd11; b = 8'd199;  #10 
a = 8'd11; b = 8'd200;  #10 
a = 8'd11; b = 8'd201;  #10 
a = 8'd11; b = 8'd202;  #10 
a = 8'd11; b = 8'd203;  #10 
a = 8'd11; b = 8'd204;  #10 
a = 8'd11; b = 8'd205;  #10 
a = 8'd11; b = 8'd206;  #10 
a = 8'd11; b = 8'd207;  #10 
a = 8'd11; b = 8'd208;  #10 
a = 8'd11; b = 8'd209;  #10 
a = 8'd11; b = 8'd210;  #10 
a = 8'd11; b = 8'd211;  #10 
a = 8'd11; b = 8'd212;  #10 
a = 8'd11; b = 8'd213;  #10 
a = 8'd11; b = 8'd214;  #10 
a = 8'd11; b = 8'd215;  #10 
a = 8'd11; b = 8'd216;  #10 
a = 8'd11; b = 8'd217;  #10 
a = 8'd11; b = 8'd218;  #10 
a = 8'd11; b = 8'd219;  #10 
a = 8'd11; b = 8'd220;  #10 
a = 8'd11; b = 8'd221;  #10 
a = 8'd11; b = 8'd222;  #10 
a = 8'd11; b = 8'd223;  #10 
a = 8'd11; b = 8'd224;  #10 
a = 8'd11; b = 8'd225;  #10 
a = 8'd11; b = 8'd226;  #10 
a = 8'd11; b = 8'd227;  #10 
a = 8'd11; b = 8'd228;  #10 
a = 8'd11; b = 8'd229;  #10 
a = 8'd11; b = 8'd230;  #10 
a = 8'd11; b = 8'd231;  #10 
a = 8'd11; b = 8'd232;  #10 
a = 8'd11; b = 8'd233;  #10 
a = 8'd11; b = 8'd234;  #10 
a = 8'd11; b = 8'd235;  #10 
a = 8'd11; b = 8'd236;  #10 
a = 8'd11; b = 8'd237;  #10 
a = 8'd11; b = 8'd238;  #10 
a = 8'd11; b = 8'd239;  #10 
a = 8'd11; b = 8'd240;  #10 
a = 8'd11; b = 8'd241;  #10 
a = 8'd11; b = 8'd242;  #10 
a = 8'd11; b = 8'd243;  #10 
a = 8'd11; b = 8'd244;  #10 
a = 8'd11; b = 8'd245;  #10 
a = 8'd11; b = 8'd246;  #10 
a = 8'd11; b = 8'd247;  #10 
a = 8'd11; b = 8'd248;  #10 
a = 8'd11; b = 8'd249;  #10 
a = 8'd11; b = 8'd250;  #10 
a = 8'd11; b = 8'd251;  #10 
a = 8'd11; b = 8'd252;  #10 
a = 8'd11; b = 8'd253;  #10 
a = 8'd11; b = 8'd254;  #10 
a = 8'd11; b = 8'd255;  #10 
a = 8'd12; b = 8'd0;  #10 
a = 8'd12; b = 8'd1;  #10 
a = 8'd12; b = 8'd2;  #10 
a = 8'd12; b = 8'd3;  #10 
a = 8'd12; b = 8'd4;  #10 
a = 8'd12; b = 8'd5;  #10 
a = 8'd12; b = 8'd6;  #10 
a = 8'd12; b = 8'd7;  #10 
a = 8'd12; b = 8'd8;  #10 
a = 8'd12; b = 8'd9;  #10 
a = 8'd12; b = 8'd10;  #10 
a = 8'd12; b = 8'd11;  #10 
a = 8'd12; b = 8'd12;  #10 
a = 8'd12; b = 8'd13;  #10 
a = 8'd12; b = 8'd14;  #10 
a = 8'd12; b = 8'd15;  #10 
a = 8'd12; b = 8'd16;  #10 
a = 8'd12; b = 8'd17;  #10 
a = 8'd12; b = 8'd18;  #10 
a = 8'd12; b = 8'd19;  #10 
a = 8'd12; b = 8'd20;  #10 
a = 8'd12; b = 8'd21;  #10 
a = 8'd12; b = 8'd22;  #10 
a = 8'd12; b = 8'd23;  #10 
a = 8'd12; b = 8'd24;  #10 
a = 8'd12; b = 8'd25;  #10 
a = 8'd12; b = 8'd26;  #10 
a = 8'd12; b = 8'd27;  #10 
a = 8'd12; b = 8'd28;  #10 
a = 8'd12; b = 8'd29;  #10 
a = 8'd12; b = 8'd30;  #10 
a = 8'd12; b = 8'd31;  #10 
a = 8'd12; b = 8'd32;  #10 
a = 8'd12; b = 8'd33;  #10 
a = 8'd12; b = 8'd34;  #10 
a = 8'd12; b = 8'd35;  #10 
a = 8'd12; b = 8'd36;  #10 
a = 8'd12; b = 8'd37;  #10 
a = 8'd12; b = 8'd38;  #10 
a = 8'd12; b = 8'd39;  #10 
a = 8'd12; b = 8'd40;  #10 
a = 8'd12; b = 8'd41;  #10 
a = 8'd12; b = 8'd42;  #10 
a = 8'd12; b = 8'd43;  #10 
a = 8'd12; b = 8'd44;  #10 
a = 8'd12; b = 8'd45;  #10 
a = 8'd12; b = 8'd46;  #10 
a = 8'd12; b = 8'd47;  #10 
a = 8'd12; b = 8'd48;  #10 
a = 8'd12; b = 8'd49;  #10 
a = 8'd12; b = 8'd50;  #10 
a = 8'd12; b = 8'd51;  #10 
a = 8'd12; b = 8'd52;  #10 
a = 8'd12; b = 8'd53;  #10 
a = 8'd12; b = 8'd54;  #10 
a = 8'd12; b = 8'd55;  #10 
a = 8'd12; b = 8'd56;  #10 
a = 8'd12; b = 8'd57;  #10 
a = 8'd12; b = 8'd58;  #10 
a = 8'd12; b = 8'd59;  #10 
a = 8'd12; b = 8'd60;  #10 
a = 8'd12; b = 8'd61;  #10 
a = 8'd12; b = 8'd62;  #10 
a = 8'd12; b = 8'd63;  #10 
a = 8'd12; b = 8'd64;  #10 
a = 8'd12; b = 8'd65;  #10 
a = 8'd12; b = 8'd66;  #10 
a = 8'd12; b = 8'd67;  #10 
a = 8'd12; b = 8'd68;  #10 
a = 8'd12; b = 8'd69;  #10 
a = 8'd12; b = 8'd70;  #10 
a = 8'd12; b = 8'd71;  #10 
a = 8'd12; b = 8'd72;  #10 
a = 8'd12; b = 8'd73;  #10 
a = 8'd12; b = 8'd74;  #10 
a = 8'd12; b = 8'd75;  #10 
a = 8'd12; b = 8'd76;  #10 
a = 8'd12; b = 8'd77;  #10 
a = 8'd12; b = 8'd78;  #10 
a = 8'd12; b = 8'd79;  #10 
a = 8'd12; b = 8'd80;  #10 
a = 8'd12; b = 8'd81;  #10 
a = 8'd12; b = 8'd82;  #10 
a = 8'd12; b = 8'd83;  #10 
a = 8'd12; b = 8'd84;  #10 
a = 8'd12; b = 8'd85;  #10 
a = 8'd12; b = 8'd86;  #10 
a = 8'd12; b = 8'd87;  #10 
a = 8'd12; b = 8'd88;  #10 
a = 8'd12; b = 8'd89;  #10 
a = 8'd12; b = 8'd90;  #10 
a = 8'd12; b = 8'd91;  #10 
a = 8'd12; b = 8'd92;  #10 
a = 8'd12; b = 8'd93;  #10 
a = 8'd12; b = 8'd94;  #10 
a = 8'd12; b = 8'd95;  #10 
a = 8'd12; b = 8'd96;  #10 
a = 8'd12; b = 8'd97;  #10 
a = 8'd12; b = 8'd98;  #10 
a = 8'd12; b = 8'd99;  #10 
a = 8'd12; b = 8'd100;  #10 
a = 8'd12; b = 8'd101;  #10 
a = 8'd12; b = 8'd102;  #10 
a = 8'd12; b = 8'd103;  #10 
a = 8'd12; b = 8'd104;  #10 
a = 8'd12; b = 8'd105;  #10 
a = 8'd12; b = 8'd106;  #10 
a = 8'd12; b = 8'd107;  #10 
a = 8'd12; b = 8'd108;  #10 
a = 8'd12; b = 8'd109;  #10 
a = 8'd12; b = 8'd110;  #10 
a = 8'd12; b = 8'd111;  #10 
a = 8'd12; b = 8'd112;  #10 
a = 8'd12; b = 8'd113;  #10 
a = 8'd12; b = 8'd114;  #10 
a = 8'd12; b = 8'd115;  #10 
a = 8'd12; b = 8'd116;  #10 
a = 8'd12; b = 8'd117;  #10 
a = 8'd12; b = 8'd118;  #10 
a = 8'd12; b = 8'd119;  #10 
a = 8'd12; b = 8'd120;  #10 
a = 8'd12; b = 8'd121;  #10 
a = 8'd12; b = 8'd122;  #10 
a = 8'd12; b = 8'd123;  #10 
a = 8'd12; b = 8'd124;  #10 
a = 8'd12; b = 8'd125;  #10 
a = 8'd12; b = 8'd126;  #10 
a = 8'd12; b = 8'd127;  #10 
a = 8'd12; b = 8'd128;  #10 
a = 8'd12; b = 8'd129;  #10 
a = 8'd12; b = 8'd130;  #10 
a = 8'd12; b = 8'd131;  #10 
a = 8'd12; b = 8'd132;  #10 
a = 8'd12; b = 8'd133;  #10 
a = 8'd12; b = 8'd134;  #10 
a = 8'd12; b = 8'd135;  #10 
a = 8'd12; b = 8'd136;  #10 
a = 8'd12; b = 8'd137;  #10 
a = 8'd12; b = 8'd138;  #10 
a = 8'd12; b = 8'd139;  #10 
a = 8'd12; b = 8'd140;  #10 
a = 8'd12; b = 8'd141;  #10 
a = 8'd12; b = 8'd142;  #10 
a = 8'd12; b = 8'd143;  #10 
a = 8'd12; b = 8'd144;  #10 
a = 8'd12; b = 8'd145;  #10 
a = 8'd12; b = 8'd146;  #10 
a = 8'd12; b = 8'd147;  #10 
a = 8'd12; b = 8'd148;  #10 
a = 8'd12; b = 8'd149;  #10 
a = 8'd12; b = 8'd150;  #10 
a = 8'd12; b = 8'd151;  #10 
a = 8'd12; b = 8'd152;  #10 
a = 8'd12; b = 8'd153;  #10 
a = 8'd12; b = 8'd154;  #10 
a = 8'd12; b = 8'd155;  #10 
a = 8'd12; b = 8'd156;  #10 
a = 8'd12; b = 8'd157;  #10 
a = 8'd12; b = 8'd158;  #10 
a = 8'd12; b = 8'd159;  #10 
a = 8'd12; b = 8'd160;  #10 
a = 8'd12; b = 8'd161;  #10 
a = 8'd12; b = 8'd162;  #10 
a = 8'd12; b = 8'd163;  #10 
a = 8'd12; b = 8'd164;  #10 
a = 8'd12; b = 8'd165;  #10 
a = 8'd12; b = 8'd166;  #10 
a = 8'd12; b = 8'd167;  #10 
a = 8'd12; b = 8'd168;  #10 
a = 8'd12; b = 8'd169;  #10 
a = 8'd12; b = 8'd170;  #10 
a = 8'd12; b = 8'd171;  #10 
a = 8'd12; b = 8'd172;  #10 
a = 8'd12; b = 8'd173;  #10 
a = 8'd12; b = 8'd174;  #10 
a = 8'd12; b = 8'd175;  #10 
a = 8'd12; b = 8'd176;  #10 
a = 8'd12; b = 8'd177;  #10 
a = 8'd12; b = 8'd178;  #10 
a = 8'd12; b = 8'd179;  #10 
a = 8'd12; b = 8'd180;  #10 
a = 8'd12; b = 8'd181;  #10 
a = 8'd12; b = 8'd182;  #10 
a = 8'd12; b = 8'd183;  #10 
a = 8'd12; b = 8'd184;  #10 
a = 8'd12; b = 8'd185;  #10 
a = 8'd12; b = 8'd186;  #10 
a = 8'd12; b = 8'd187;  #10 
a = 8'd12; b = 8'd188;  #10 
a = 8'd12; b = 8'd189;  #10 
a = 8'd12; b = 8'd190;  #10 
a = 8'd12; b = 8'd191;  #10 
a = 8'd12; b = 8'd192;  #10 
a = 8'd12; b = 8'd193;  #10 
a = 8'd12; b = 8'd194;  #10 
a = 8'd12; b = 8'd195;  #10 
a = 8'd12; b = 8'd196;  #10 
a = 8'd12; b = 8'd197;  #10 
a = 8'd12; b = 8'd198;  #10 
a = 8'd12; b = 8'd199;  #10 
a = 8'd12; b = 8'd200;  #10 
a = 8'd12; b = 8'd201;  #10 
a = 8'd12; b = 8'd202;  #10 
a = 8'd12; b = 8'd203;  #10 
a = 8'd12; b = 8'd204;  #10 
a = 8'd12; b = 8'd205;  #10 
a = 8'd12; b = 8'd206;  #10 
a = 8'd12; b = 8'd207;  #10 
a = 8'd12; b = 8'd208;  #10 
a = 8'd12; b = 8'd209;  #10 
a = 8'd12; b = 8'd210;  #10 
a = 8'd12; b = 8'd211;  #10 
a = 8'd12; b = 8'd212;  #10 
a = 8'd12; b = 8'd213;  #10 
a = 8'd12; b = 8'd214;  #10 
a = 8'd12; b = 8'd215;  #10 
a = 8'd12; b = 8'd216;  #10 
a = 8'd12; b = 8'd217;  #10 
a = 8'd12; b = 8'd218;  #10 
a = 8'd12; b = 8'd219;  #10 
a = 8'd12; b = 8'd220;  #10 
a = 8'd12; b = 8'd221;  #10 
a = 8'd12; b = 8'd222;  #10 
a = 8'd12; b = 8'd223;  #10 
a = 8'd12; b = 8'd224;  #10 
a = 8'd12; b = 8'd225;  #10 
a = 8'd12; b = 8'd226;  #10 
a = 8'd12; b = 8'd227;  #10 
a = 8'd12; b = 8'd228;  #10 
a = 8'd12; b = 8'd229;  #10 
a = 8'd12; b = 8'd230;  #10 
a = 8'd12; b = 8'd231;  #10 
a = 8'd12; b = 8'd232;  #10 
a = 8'd12; b = 8'd233;  #10 
a = 8'd12; b = 8'd234;  #10 
a = 8'd12; b = 8'd235;  #10 
a = 8'd12; b = 8'd236;  #10 
a = 8'd12; b = 8'd237;  #10 
a = 8'd12; b = 8'd238;  #10 
a = 8'd12; b = 8'd239;  #10 
a = 8'd12; b = 8'd240;  #10 
a = 8'd12; b = 8'd241;  #10 
a = 8'd12; b = 8'd242;  #10 
a = 8'd12; b = 8'd243;  #10 
a = 8'd12; b = 8'd244;  #10 
a = 8'd12; b = 8'd245;  #10 
a = 8'd12; b = 8'd246;  #10 
a = 8'd12; b = 8'd247;  #10 
a = 8'd12; b = 8'd248;  #10 
a = 8'd12; b = 8'd249;  #10 
a = 8'd12; b = 8'd250;  #10 
a = 8'd12; b = 8'd251;  #10 
a = 8'd12; b = 8'd252;  #10 
a = 8'd12; b = 8'd253;  #10 
a = 8'd12; b = 8'd254;  #10 
a = 8'd12; b = 8'd255;  #10 
a = 8'd13; b = 8'd0;  #10 
a = 8'd13; b = 8'd1;  #10 
a = 8'd13; b = 8'd2;  #10 
a = 8'd13; b = 8'd3;  #10 
a = 8'd13; b = 8'd4;  #10 
a = 8'd13; b = 8'd5;  #10 
a = 8'd13; b = 8'd6;  #10 
a = 8'd13; b = 8'd7;  #10 
a = 8'd13; b = 8'd8;  #10 
a = 8'd13; b = 8'd9;  #10 
a = 8'd13; b = 8'd10;  #10 
a = 8'd13; b = 8'd11;  #10 
a = 8'd13; b = 8'd12;  #10 
a = 8'd13; b = 8'd13;  #10 
a = 8'd13; b = 8'd14;  #10 
a = 8'd13; b = 8'd15;  #10 
a = 8'd13; b = 8'd16;  #10 
a = 8'd13; b = 8'd17;  #10 
a = 8'd13; b = 8'd18;  #10 
a = 8'd13; b = 8'd19;  #10 
a = 8'd13; b = 8'd20;  #10 
a = 8'd13; b = 8'd21;  #10 
a = 8'd13; b = 8'd22;  #10 
a = 8'd13; b = 8'd23;  #10 
a = 8'd13; b = 8'd24;  #10 
a = 8'd13; b = 8'd25;  #10 
a = 8'd13; b = 8'd26;  #10 
a = 8'd13; b = 8'd27;  #10 
a = 8'd13; b = 8'd28;  #10 
a = 8'd13; b = 8'd29;  #10 
a = 8'd13; b = 8'd30;  #10 
a = 8'd13; b = 8'd31;  #10 
a = 8'd13; b = 8'd32;  #10 
a = 8'd13; b = 8'd33;  #10 
a = 8'd13; b = 8'd34;  #10 
a = 8'd13; b = 8'd35;  #10 
a = 8'd13; b = 8'd36;  #10 
a = 8'd13; b = 8'd37;  #10 
a = 8'd13; b = 8'd38;  #10 
a = 8'd13; b = 8'd39;  #10 
a = 8'd13; b = 8'd40;  #10 
a = 8'd13; b = 8'd41;  #10 
a = 8'd13; b = 8'd42;  #10 
a = 8'd13; b = 8'd43;  #10 
a = 8'd13; b = 8'd44;  #10 
a = 8'd13; b = 8'd45;  #10 
a = 8'd13; b = 8'd46;  #10 
a = 8'd13; b = 8'd47;  #10 
a = 8'd13; b = 8'd48;  #10 
a = 8'd13; b = 8'd49;  #10 
a = 8'd13; b = 8'd50;  #10 
a = 8'd13; b = 8'd51;  #10 
a = 8'd13; b = 8'd52;  #10 
a = 8'd13; b = 8'd53;  #10 
a = 8'd13; b = 8'd54;  #10 
a = 8'd13; b = 8'd55;  #10 
a = 8'd13; b = 8'd56;  #10 
a = 8'd13; b = 8'd57;  #10 
a = 8'd13; b = 8'd58;  #10 
a = 8'd13; b = 8'd59;  #10 
a = 8'd13; b = 8'd60;  #10 
a = 8'd13; b = 8'd61;  #10 
a = 8'd13; b = 8'd62;  #10 
a = 8'd13; b = 8'd63;  #10 
a = 8'd13; b = 8'd64;  #10 
a = 8'd13; b = 8'd65;  #10 
a = 8'd13; b = 8'd66;  #10 
a = 8'd13; b = 8'd67;  #10 
a = 8'd13; b = 8'd68;  #10 
a = 8'd13; b = 8'd69;  #10 
a = 8'd13; b = 8'd70;  #10 
a = 8'd13; b = 8'd71;  #10 
a = 8'd13; b = 8'd72;  #10 
a = 8'd13; b = 8'd73;  #10 
a = 8'd13; b = 8'd74;  #10 
a = 8'd13; b = 8'd75;  #10 
a = 8'd13; b = 8'd76;  #10 
a = 8'd13; b = 8'd77;  #10 
a = 8'd13; b = 8'd78;  #10 
a = 8'd13; b = 8'd79;  #10 
a = 8'd13; b = 8'd80;  #10 
a = 8'd13; b = 8'd81;  #10 
a = 8'd13; b = 8'd82;  #10 
a = 8'd13; b = 8'd83;  #10 
a = 8'd13; b = 8'd84;  #10 
a = 8'd13; b = 8'd85;  #10 
a = 8'd13; b = 8'd86;  #10 
a = 8'd13; b = 8'd87;  #10 
a = 8'd13; b = 8'd88;  #10 
a = 8'd13; b = 8'd89;  #10 
a = 8'd13; b = 8'd90;  #10 
a = 8'd13; b = 8'd91;  #10 
a = 8'd13; b = 8'd92;  #10 
a = 8'd13; b = 8'd93;  #10 
a = 8'd13; b = 8'd94;  #10 
a = 8'd13; b = 8'd95;  #10 
a = 8'd13; b = 8'd96;  #10 
a = 8'd13; b = 8'd97;  #10 
a = 8'd13; b = 8'd98;  #10 
a = 8'd13; b = 8'd99;  #10 
a = 8'd13; b = 8'd100;  #10 
a = 8'd13; b = 8'd101;  #10 
a = 8'd13; b = 8'd102;  #10 
a = 8'd13; b = 8'd103;  #10 
a = 8'd13; b = 8'd104;  #10 
a = 8'd13; b = 8'd105;  #10 
a = 8'd13; b = 8'd106;  #10 
a = 8'd13; b = 8'd107;  #10 
a = 8'd13; b = 8'd108;  #10 
a = 8'd13; b = 8'd109;  #10 
a = 8'd13; b = 8'd110;  #10 
a = 8'd13; b = 8'd111;  #10 
a = 8'd13; b = 8'd112;  #10 
a = 8'd13; b = 8'd113;  #10 
a = 8'd13; b = 8'd114;  #10 
a = 8'd13; b = 8'd115;  #10 
a = 8'd13; b = 8'd116;  #10 
a = 8'd13; b = 8'd117;  #10 
a = 8'd13; b = 8'd118;  #10 
a = 8'd13; b = 8'd119;  #10 
a = 8'd13; b = 8'd120;  #10 
a = 8'd13; b = 8'd121;  #10 
a = 8'd13; b = 8'd122;  #10 
a = 8'd13; b = 8'd123;  #10 
a = 8'd13; b = 8'd124;  #10 
a = 8'd13; b = 8'd125;  #10 
a = 8'd13; b = 8'd126;  #10 
a = 8'd13; b = 8'd127;  #10 
a = 8'd13; b = 8'd128;  #10 
a = 8'd13; b = 8'd129;  #10 
a = 8'd13; b = 8'd130;  #10 
a = 8'd13; b = 8'd131;  #10 
a = 8'd13; b = 8'd132;  #10 
a = 8'd13; b = 8'd133;  #10 
a = 8'd13; b = 8'd134;  #10 
a = 8'd13; b = 8'd135;  #10 
a = 8'd13; b = 8'd136;  #10 
a = 8'd13; b = 8'd137;  #10 
a = 8'd13; b = 8'd138;  #10 
a = 8'd13; b = 8'd139;  #10 
a = 8'd13; b = 8'd140;  #10 
a = 8'd13; b = 8'd141;  #10 
a = 8'd13; b = 8'd142;  #10 
a = 8'd13; b = 8'd143;  #10 
a = 8'd13; b = 8'd144;  #10 
a = 8'd13; b = 8'd145;  #10 
a = 8'd13; b = 8'd146;  #10 
a = 8'd13; b = 8'd147;  #10 
a = 8'd13; b = 8'd148;  #10 
a = 8'd13; b = 8'd149;  #10 
a = 8'd13; b = 8'd150;  #10 
a = 8'd13; b = 8'd151;  #10 
a = 8'd13; b = 8'd152;  #10 
a = 8'd13; b = 8'd153;  #10 
a = 8'd13; b = 8'd154;  #10 
a = 8'd13; b = 8'd155;  #10 
a = 8'd13; b = 8'd156;  #10 
a = 8'd13; b = 8'd157;  #10 
a = 8'd13; b = 8'd158;  #10 
a = 8'd13; b = 8'd159;  #10 
a = 8'd13; b = 8'd160;  #10 
a = 8'd13; b = 8'd161;  #10 
a = 8'd13; b = 8'd162;  #10 
a = 8'd13; b = 8'd163;  #10 
a = 8'd13; b = 8'd164;  #10 
a = 8'd13; b = 8'd165;  #10 
a = 8'd13; b = 8'd166;  #10 
a = 8'd13; b = 8'd167;  #10 
a = 8'd13; b = 8'd168;  #10 
a = 8'd13; b = 8'd169;  #10 
a = 8'd13; b = 8'd170;  #10 
a = 8'd13; b = 8'd171;  #10 
a = 8'd13; b = 8'd172;  #10 
a = 8'd13; b = 8'd173;  #10 
a = 8'd13; b = 8'd174;  #10 
a = 8'd13; b = 8'd175;  #10 
a = 8'd13; b = 8'd176;  #10 
a = 8'd13; b = 8'd177;  #10 
a = 8'd13; b = 8'd178;  #10 
a = 8'd13; b = 8'd179;  #10 
a = 8'd13; b = 8'd180;  #10 
a = 8'd13; b = 8'd181;  #10 
a = 8'd13; b = 8'd182;  #10 
a = 8'd13; b = 8'd183;  #10 
a = 8'd13; b = 8'd184;  #10 
a = 8'd13; b = 8'd185;  #10 
a = 8'd13; b = 8'd186;  #10 
a = 8'd13; b = 8'd187;  #10 
a = 8'd13; b = 8'd188;  #10 
a = 8'd13; b = 8'd189;  #10 
a = 8'd13; b = 8'd190;  #10 
a = 8'd13; b = 8'd191;  #10 
a = 8'd13; b = 8'd192;  #10 
a = 8'd13; b = 8'd193;  #10 
a = 8'd13; b = 8'd194;  #10 
a = 8'd13; b = 8'd195;  #10 
a = 8'd13; b = 8'd196;  #10 
a = 8'd13; b = 8'd197;  #10 
a = 8'd13; b = 8'd198;  #10 
a = 8'd13; b = 8'd199;  #10 
a = 8'd13; b = 8'd200;  #10 
a = 8'd13; b = 8'd201;  #10 
a = 8'd13; b = 8'd202;  #10 
a = 8'd13; b = 8'd203;  #10 
a = 8'd13; b = 8'd204;  #10 
a = 8'd13; b = 8'd205;  #10 
a = 8'd13; b = 8'd206;  #10 
a = 8'd13; b = 8'd207;  #10 
a = 8'd13; b = 8'd208;  #10 
a = 8'd13; b = 8'd209;  #10 
a = 8'd13; b = 8'd210;  #10 
a = 8'd13; b = 8'd211;  #10 
a = 8'd13; b = 8'd212;  #10 
a = 8'd13; b = 8'd213;  #10 
a = 8'd13; b = 8'd214;  #10 
a = 8'd13; b = 8'd215;  #10 
a = 8'd13; b = 8'd216;  #10 
a = 8'd13; b = 8'd217;  #10 
a = 8'd13; b = 8'd218;  #10 
a = 8'd13; b = 8'd219;  #10 
a = 8'd13; b = 8'd220;  #10 
a = 8'd13; b = 8'd221;  #10 
a = 8'd13; b = 8'd222;  #10 
a = 8'd13; b = 8'd223;  #10 
a = 8'd13; b = 8'd224;  #10 
a = 8'd13; b = 8'd225;  #10 
a = 8'd13; b = 8'd226;  #10 
a = 8'd13; b = 8'd227;  #10 
a = 8'd13; b = 8'd228;  #10 
a = 8'd13; b = 8'd229;  #10 
a = 8'd13; b = 8'd230;  #10 
a = 8'd13; b = 8'd231;  #10 
a = 8'd13; b = 8'd232;  #10 
a = 8'd13; b = 8'd233;  #10 
a = 8'd13; b = 8'd234;  #10 
a = 8'd13; b = 8'd235;  #10 
a = 8'd13; b = 8'd236;  #10 
a = 8'd13; b = 8'd237;  #10 
a = 8'd13; b = 8'd238;  #10 
a = 8'd13; b = 8'd239;  #10 
a = 8'd13; b = 8'd240;  #10 
a = 8'd13; b = 8'd241;  #10 
a = 8'd13; b = 8'd242;  #10 
a = 8'd13; b = 8'd243;  #10 
a = 8'd13; b = 8'd244;  #10 
a = 8'd13; b = 8'd245;  #10 
a = 8'd13; b = 8'd246;  #10 
a = 8'd13; b = 8'd247;  #10 
a = 8'd13; b = 8'd248;  #10 
a = 8'd13; b = 8'd249;  #10 
a = 8'd13; b = 8'd250;  #10 
a = 8'd13; b = 8'd251;  #10 
a = 8'd13; b = 8'd252;  #10 
a = 8'd13; b = 8'd253;  #10 
a = 8'd13; b = 8'd254;  #10 
a = 8'd13; b = 8'd255;  #10 
a = 8'd14; b = 8'd0;  #10 
a = 8'd14; b = 8'd1;  #10 
a = 8'd14; b = 8'd2;  #10 
a = 8'd14; b = 8'd3;  #10 
a = 8'd14; b = 8'd4;  #10 
a = 8'd14; b = 8'd5;  #10 
a = 8'd14; b = 8'd6;  #10 
a = 8'd14; b = 8'd7;  #10 
a = 8'd14; b = 8'd8;  #10 
a = 8'd14; b = 8'd9;  #10 
a = 8'd14; b = 8'd10;  #10 
a = 8'd14; b = 8'd11;  #10 
a = 8'd14; b = 8'd12;  #10 
a = 8'd14; b = 8'd13;  #10 
a = 8'd14; b = 8'd14;  #10 
a = 8'd14; b = 8'd15;  #10 
a = 8'd14; b = 8'd16;  #10 
a = 8'd14; b = 8'd17;  #10 
a = 8'd14; b = 8'd18;  #10 
a = 8'd14; b = 8'd19;  #10 
a = 8'd14; b = 8'd20;  #10 
a = 8'd14; b = 8'd21;  #10 
a = 8'd14; b = 8'd22;  #10 
a = 8'd14; b = 8'd23;  #10 
a = 8'd14; b = 8'd24;  #10 
a = 8'd14; b = 8'd25;  #10 
a = 8'd14; b = 8'd26;  #10 
a = 8'd14; b = 8'd27;  #10 
a = 8'd14; b = 8'd28;  #10 
a = 8'd14; b = 8'd29;  #10 
a = 8'd14; b = 8'd30;  #10 
a = 8'd14; b = 8'd31;  #10 
a = 8'd14; b = 8'd32;  #10 
a = 8'd14; b = 8'd33;  #10 
a = 8'd14; b = 8'd34;  #10 
a = 8'd14; b = 8'd35;  #10 
a = 8'd14; b = 8'd36;  #10 
a = 8'd14; b = 8'd37;  #10 
a = 8'd14; b = 8'd38;  #10 
a = 8'd14; b = 8'd39;  #10 
a = 8'd14; b = 8'd40;  #10 
a = 8'd14; b = 8'd41;  #10 
a = 8'd14; b = 8'd42;  #10 
a = 8'd14; b = 8'd43;  #10 
a = 8'd14; b = 8'd44;  #10 
a = 8'd14; b = 8'd45;  #10 
a = 8'd14; b = 8'd46;  #10 
a = 8'd14; b = 8'd47;  #10 
a = 8'd14; b = 8'd48;  #10 
a = 8'd14; b = 8'd49;  #10 
a = 8'd14; b = 8'd50;  #10 
a = 8'd14; b = 8'd51;  #10 
a = 8'd14; b = 8'd52;  #10 
a = 8'd14; b = 8'd53;  #10 
a = 8'd14; b = 8'd54;  #10 
a = 8'd14; b = 8'd55;  #10 
a = 8'd14; b = 8'd56;  #10 
a = 8'd14; b = 8'd57;  #10 
a = 8'd14; b = 8'd58;  #10 
a = 8'd14; b = 8'd59;  #10 
a = 8'd14; b = 8'd60;  #10 
a = 8'd14; b = 8'd61;  #10 
a = 8'd14; b = 8'd62;  #10 
a = 8'd14; b = 8'd63;  #10 
a = 8'd14; b = 8'd64;  #10 
a = 8'd14; b = 8'd65;  #10 
a = 8'd14; b = 8'd66;  #10 
a = 8'd14; b = 8'd67;  #10 
a = 8'd14; b = 8'd68;  #10 
a = 8'd14; b = 8'd69;  #10 
a = 8'd14; b = 8'd70;  #10 
a = 8'd14; b = 8'd71;  #10 
a = 8'd14; b = 8'd72;  #10 
a = 8'd14; b = 8'd73;  #10 
a = 8'd14; b = 8'd74;  #10 
a = 8'd14; b = 8'd75;  #10 
a = 8'd14; b = 8'd76;  #10 
a = 8'd14; b = 8'd77;  #10 
a = 8'd14; b = 8'd78;  #10 
a = 8'd14; b = 8'd79;  #10 
a = 8'd14; b = 8'd80;  #10 
a = 8'd14; b = 8'd81;  #10 
a = 8'd14; b = 8'd82;  #10 
a = 8'd14; b = 8'd83;  #10 
a = 8'd14; b = 8'd84;  #10 
a = 8'd14; b = 8'd85;  #10 
a = 8'd14; b = 8'd86;  #10 
a = 8'd14; b = 8'd87;  #10 
a = 8'd14; b = 8'd88;  #10 
a = 8'd14; b = 8'd89;  #10 
a = 8'd14; b = 8'd90;  #10 
a = 8'd14; b = 8'd91;  #10 
a = 8'd14; b = 8'd92;  #10 
a = 8'd14; b = 8'd93;  #10 
a = 8'd14; b = 8'd94;  #10 
a = 8'd14; b = 8'd95;  #10 
a = 8'd14; b = 8'd96;  #10 
a = 8'd14; b = 8'd97;  #10 
a = 8'd14; b = 8'd98;  #10 
a = 8'd14; b = 8'd99;  #10 
a = 8'd14; b = 8'd100;  #10 
a = 8'd14; b = 8'd101;  #10 
a = 8'd14; b = 8'd102;  #10 
a = 8'd14; b = 8'd103;  #10 
a = 8'd14; b = 8'd104;  #10 
a = 8'd14; b = 8'd105;  #10 
a = 8'd14; b = 8'd106;  #10 
a = 8'd14; b = 8'd107;  #10 
a = 8'd14; b = 8'd108;  #10 
a = 8'd14; b = 8'd109;  #10 
a = 8'd14; b = 8'd110;  #10 
a = 8'd14; b = 8'd111;  #10 
a = 8'd14; b = 8'd112;  #10 
a = 8'd14; b = 8'd113;  #10 
a = 8'd14; b = 8'd114;  #10 
a = 8'd14; b = 8'd115;  #10 
a = 8'd14; b = 8'd116;  #10 
a = 8'd14; b = 8'd117;  #10 
a = 8'd14; b = 8'd118;  #10 
a = 8'd14; b = 8'd119;  #10 
a = 8'd14; b = 8'd120;  #10 
a = 8'd14; b = 8'd121;  #10 
a = 8'd14; b = 8'd122;  #10 
a = 8'd14; b = 8'd123;  #10 
a = 8'd14; b = 8'd124;  #10 
a = 8'd14; b = 8'd125;  #10 
a = 8'd14; b = 8'd126;  #10 
a = 8'd14; b = 8'd127;  #10 
a = 8'd14; b = 8'd128;  #10 
a = 8'd14; b = 8'd129;  #10 
a = 8'd14; b = 8'd130;  #10 
a = 8'd14; b = 8'd131;  #10 
a = 8'd14; b = 8'd132;  #10 
a = 8'd14; b = 8'd133;  #10 
a = 8'd14; b = 8'd134;  #10 
a = 8'd14; b = 8'd135;  #10 
a = 8'd14; b = 8'd136;  #10 
a = 8'd14; b = 8'd137;  #10 
a = 8'd14; b = 8'd138;  #10 
a = 8'd14; b = 8'd139;  #10 
a = 8'd14; b = 8'd140;  #10 
a = 8'd14; b = 8'd141;  #10 
a = 8'd14; b = 8'd142;  #10 
a = 8'd14; b = 8'd143;  #10 
a = 8'd14; b = 8'd144;  #10 
a = 8'd14; b = 8'd145;  #10 
a = 8'd14; b = 8'd146;  #10 
a = 8'd14; b = 8'd147;  #10 
a = 8'd14; b = 8'd148;  #10 
a = 8'd14; b = 8'd149;  #10 
a = 8'd14; b = 8'd150;  #10 
a = 8'd14; b = 8'd151;  #10 
a = 8'd14; b = 8'd152;  #10 
a = 8'd14; b = 8'd153;  #10 
a = 8'd14; b = 8'd154;  #10 
a = 8'd14; b = 8'd155;  #10 
a = 8'd14; b = 8'd156;  #10 
a = 8'd14; b = 8'd157;  #10 
a = 8'd14; b = 8'd158;  #10 
a = 8'd14; b = 8'd159;  #10 
a = 8'd14; b = 8'd160;  #10 
a = 8'd14; b = 8'd161;  #10 
a = 8'd14; b = 8'd162;  #10 
a = 8'd14; b = 8'd163;  #10 
a = 8'd14; b = 8'd164;  #10 
a = 8'd14; b = 8'd165;  #10 
a = 8'd14; b = 8'd166;  #10 
a = 8'd14; b = 8'd167;  #10 
a = 8'd14; b = 8'd168;  #10 
a = 8'd14; b = 8'd169;  #10 
a = 8'd14; b = 8'd170;  #10 
a = 8'd14; b = 8'd171;  #10 
a = 8'd14; b = 8'd172;  #10 
a = 8'd14; b = 8'd173;  #10 
a = 8'd14; b = 8'd174;  #10 
a = 8'd14; b = 8'd175;  #10 
a = 8'd14; b = 8'd176;  #10 
a = 8'd14; b = 8'd177;  #10 
a = 8'd14; b = 8'd178;  #10 
a = 8'd14; b = 8'd179;  #10 
a = 8'd14; b = 8'd180;  #10 
a = 8'd14; b = 8'd181;  #10 
a = 8'd14; b = 8'd182;  #10 
a = 8'd14; b = 8'd183;  #10 
a = 8'd14; b = 8'd184;  #10 
a = 8'd14; b = 8'd185;  #10 
a = 8'd14; b = 8'd186;  #10 
a = 8'd14; b = 8'd187;  #10 
a = 8'd14; b = 8'd188;  #10 
a = 8'd14; b = 8'd189;  #10 
a = 8'd14; b = 8'd190;  #10 
a = 8'd14; b = 8'd191;  #10 
a = 8'd14; b = 8'd192;  #10 
a = 8'd14; b = 8'd193;  #10 
a = 8'd14; b = 8'd194;  #10 
a = 8'd14; b = 8'd195;  #10 
a = 8'd14; b = 8'd196;  #10 
a = 8'd14; b = 8'd197;  #10 
a = 8'd14; b = 8'd198;  #10 
a = 8'd14; b = 8'd199;  #10 
a = 8'd14; b = 8'd200;  #10 
a = 8'd14; b = 8'd201;  #10 
a = 8'd14; b = 8'd202;  #10 
a = 8'd14; b = 8'd203;  #10 
a = 8'd14; b = 8'd204;  #10 
a = 8'd14; b = 8'd205;  #10 
a = 8'd14; b = 8'd206;  #10 
a = 8'd14; b = 8'd207;  #10 
a = 8'd14; b = 8'd208;  #10 
a = 8'd14; b = 8'd209;  #10 
a = 8'd14; b = 8'd210;  #10 
a = 8'd14; b = 8'd211;  #10 
a = 8'd14; b = 8'd212;  #10 
a = 8'd14; b = 8'd213;  #10 
a = 8'd14; b = 8'd214;  #10 
a = 8'd14; b = 8'd215;  #10 
a = 8'd14; b = 8'd216;  #10 
a = 8'd14; b = 8'd217;  #10 
a = 8'd14; b = 8'd218;  #10 
a = 8'd14; b = 8'd219;  #10 
a = 8'd14; b = 8'd220;  #10 
a = 8'd14; b = 8'd221;  #10 
a = 8'd14; b = 8'd222;  #10 
a = 8'd14; b = 8'd223;  #10 
a = 8'd14; b = 8'd224;  #10 
a = 8'd14; b = 8'd225;  #10 
a = 8'd14; b = 8'd226;  #10 
a = 8'd14; b = 8'd227;  #10 
a = 8'd14; b = 8'd228;  #10 
a = 8'd14; b = 8'd229;  #10 
a = 8'd14; b = 8'd230;  #10 
a = 8'd14; b = 8'd231;  #10 
a = 8'd14; b = 8'd232;  #10 
a = 8'd14; b = 8'd233;  #10 
a = 8'd14; b = 8'd234;  #10 
a = 8'd14; b = 8'd235;  #10 
a = 8'd14; b = 8'd236;  #10 
a = 8'd14; b = 8'd237;  #10 
a = 8'd14; b = 8'd238;  #10 
a = 8'd14; b = 8'd239;  #10 
a = 8'd14; b = 8'd240;  #10 
a = 8'd14; b = 8'd241;  #10 
a = 8'd14; b = 8'd242;  #10 
a = 8'd14; b = 8'd243;  #10 
a = 8'd14; b = 8'd244;  #10 
a = 8'd14; b = 8'd245;  #10 
a = 8'd14; b = 8'd246;  #10 
a = 8'd14; b = 8'd247;  #10 
a = 8'd14; b = 8'd248;  #10 
a = 8'd14; b = 8'd249;  #10 
a = 8'd14; b = 8'd250;  #10 
a = 8'd14; b = 8'd251;  #10 
a = 8'd14; b = 8'd252;  #10 
a = 8'd14; b = 8'd253;  #10 
a = 8'd14; b = 8'd254;  #10 
a = 8'd14; b = 8'd255;  #10 
a = 8'd15; b = 8'd0;  #10 
a = 8'd15; b = 8'd1;  #10 
a = 8'd15; b = 8'd2;  #10 
a = 8'd15; b = 8'd3;  #10 
a = 8'd15; b = 8'd4;  #10 
a = 8'd15; b = 8'd5;  #10 
a = 8'd15; b = 8'd6;  #10 
a = 8'd15; b = 8'd7;  #10 
a = 8'd15; b = 8'd8;  #10 
a = 8'd15; b = 8'd9;  #10 
a = 8'd15; b = 8'd10;  #10 
a = 8'd15; b = 8'd11;  #10 
a = 8'd15; b = 8'd12;  #10 
a = 8'd15; b = 8'd13;  #10 
a = 8'd15; b = 8'd14;  #10 
a = 8'd15; b = 8'd15;  #10 
a = 8'd15; b = 8'd16;  #10 
a = 8'd15; b = 8'd17;  #10 
a = 8'd15; b = 8'd18;  #10 
a = 8'd15; b = 8'd19;  #10 
a = 8'd15; b = 8'd20;  #10 
a = 8'd15; b = 8'd21;  #10 
a = 8'd15; b = 8'd22;  #10 
a = 8'd15; b = 8'd23;  #10 
a = 8'd15; b = 8'd24;  #10 
a = 8'd15; b = 8'd25;  #10 
a = 8'd15; b = 8'd26;  #10 
a = 8'd15; b = 8'd27;  #10 
a = 8'd15; b = 8'd28;  #10 
a = 8'd15; b = 8'd29;  #10 
a = 8'd15; b = 8'd30;  #10 
a = 8'd15; b = 8'd31;  #10 
a = 8'd15; b = 8'd32;  #10 
a = 8'd15; b = 8'd33;  #10 
a = 8'd15; b = 8'd34;  #10 
a = 8'd15; b = 8'd35;  #10 
a = 8'd15; b = 8'd36;  #10 
a = 8'd15; b = 8'd37;  #10 
a = 8'd15; b = 8'd38;  #10 
a = 8'd15; b = 8'd39;  #10 
a = 8'd15; b = 8'd40;  #10 
a = 8'd15; b = 8'd41;  #10 
a = 8'd15; b = 8'd42;  #10 
a = 8'd15; b = 8'd43;  #10 
a = 8'd15; b = 8'd44;  #10 
a = 8'd15; b = 8'd45;  #10 
a = 8'd15; b = 8'd46;  #10 
a = 8'd15; b = 8'd47;  #10 
a = 8'd15; b = 8'd48;  #10 
a = 8'd15; b = 8'd49;  #10 
a = 8'd15; b = 8'd50;  #10 
a = 8'd15; b = 8'd51;  #10 
a = 8'd15; b = 8'd52;  #10 
a = 8'd15; b = 8'd53;  #10 
a = 8'd15; b = 8'd54;  #10 
a = 8'd15; b = 8'd55;  #10 
a = 8'd15; b = 8'd56;  #10 
a = 8'd15; b = 8'd57;  #10 
a = 8'd15; b = 8'd58;  #10 
a = 8'd15; b = 8'd59;  #10 
a = 8'd15; b = 8'd60;  #10 
a = 8'd15; b = 8'd61;  #10 
a = 8'd15; b = 8'd62;  #10 
a = 8'd15; b = 8'd63;  #10 
a = 8'd15; b = 8'd64;  #10 
a = 8'd15; b = 8'd65;  #10 
a = 8'd15; b = 8'd66;  #10 
a = 8'd15; b = 8'd67;  #10 
a = 8'd15; b = 8'd68;  #10 
a = 8'd15; b = 8'd69;  #10 
a = 8'd15; b = 8'd70;  #10 
a = 8'd15; b = 8'd71;  #10 
a = 8'd15; b = 8'd72;  #10 
a = 8'd15; b = 8'd73;  #10 
a = 8'd15; b = 8'd74;  #10 
a = 8'd15; b = 8'd75;  #10 
a = 8'd15; b = 8'd76;  #10 
a = 8'd15; b = 8'd77;  #10 
a = 8'd15; b = 8'd78;  #10 
a = 8'd15; b = 8'd79;  #10 
a = 8'd15; b = 8'd80;  #10 
a = 8'd15; b = 8'd81;  #10 
a = 8'd15; b = 8'd82;  #10 
a = 8'd15; b = 8'd83;  #10 
a = 8'd15; b = 8'd84;  #10 
a = 8'd15; b = 8'd85;  #10 
a = 8'd15; b = 8'd86;  #10 
a = 8'd15; b = 8'd87;  #10 
a = 8'd15; b = 8'd88;  #10 
a = 8'd15; b = 8'd89;  #10 
a = 8'd15; b = 8'd90;  #10 
a = 8'd15; b = 8'd91;  #10 
a = 8'd15; b = 8'd92;  #10 
a = 8'd15; b = 8'd93;  #10 
a = 8'd15; b = 8'd94;  #10 
a = 8'd15; b = 8'd95;  #10 
a = 8'd15; b = 8'd96;  #10 
a = 8'd15; b = 8'd97;  #10 
a = 8'd15; b = 8'd98;  #10 
a = 8'd15; b = 8'd99;  #10 
a = 8'd15; b = 8'd100;  #10 
a = 8'd15; b = 8'd101;  #10 
a = 8'd15; b = 8'd102;  #10 
a = 8'd15; b = 8'd103;  #10 
a = 8'd15; b = 8'd104;  #10 
a = 8'd15; b = 8'd105;  #10 
a = 8'd15; b = 8'd106;  #10 
a = 8'd15; b = 8'd107;  #10 
a = 8'd15; b = 8'd108;  #10 
a = 8'd15; b = 8'd109;  #10 
a = 8'd15; b = 8'd110;  #10 
a = 8'd15; b = 8'd111;  #10 
a = 8'd15; b = 8'd112;  #10 
a = 8'd15; b = 8'd113;  #10 
a = 8'd15; b = 8'd114;  #10 
a = 8'd15; b = 8'd115;  #10 
a = 8'd15; b = 8'd116;  #10 
a = 8'd15; b = 8'd117;  #10 
a = 8'd15; b = 8'd118;  #10 
a = 8'd15; b = 8'd119;  #10 
a = 8'd15; b = 8'd120;  #10 
a = 8'd15; b = 8'd121;  #10 
a = 8'd15; b = 8'd122;  #10 
a = 8'd15; b = 8'd123;  #10 
a = 8'd15; b = 8'd124;  #10 
a = 8'd15; b = 8'd125;  #10 
a = 8'd15; b = 8'd126;  #10 
a = 8'd15; b = 8'd127;  #10 
a = 8'd15; b = 8'd128;  #10 
a = 8'd15; b = 8'd129;  #10 
a = 8'd15; b = 8'd130;  #10 
a = 8'd15; b = 8'd131;  #10 
a = 8'd15; b = 8'd132;  #10 
a = 8'd15; b = 8'd133;  #10 
a = 8'd15; b = 8'd134;  #10 
a = 8'd15; b = 8'd135;  #10 
a = 8'd15; b = 8'd136;  #10 
a = 8'd15; b = 8'd137;  #10 
a = 8'd15; b = 8'd138;  #10 
a = 8'd15; b = 8'd139;  #10 
a = 8'd15; b = 8'd140;  #10 
a = 8'd15; b = 8'd141;  #10 
a = 8'd15; b = 8'd142;  #10 
a = 8'd15; b = 8'd143;  #10 
a = 8'd15; b = 8'd144;  #10 
a = 8'd15; b = 8'd145;  #10 
a = 8'd15; b = 8'd146;  #10 
a = 8'd15; b = 8'd147;  #10 
a = 8'd15; b = 8'd148;  #10 
a = 8'd15; b = 8'd149;  #10 
a = 8'd15; b = 8'd150;  #10 
a = 8'd15; b = 8'd151;  #10 
a = 8'd15; b = 8'd152;  #10 
a = 8'd15; b = 8'd153;  #10 
a = 8'd15; b = 8'd154;  #10 
a = 8'd15; b = 8'd155;  #10 
a = 8'd15; b = 8'd156;  #10 
a = 8'd15; b = 8'd157;  #10 
a = 8'd15; b = 8'd158;  #10 
a = 8'd15; b = 8'd159;  #10 
a = 8'd15; b = 8'd160;  #10 
a = 8'd15; b = 8'd161;  #10 
a = 8'd15; b = 8'd162;  #10 
a = 8'd15; b = 8'd163;  #10 
a = 8'd15; b = 8'd164;  #10 
a = 8'd15; b = 8'd165;  #10 
a = 8'd15; b = 8'd166;  #10 
a = 8'd15; b = 8'd167;  #10 
a = 8'd15; b = 8'd168;  #10 
a = 8'd15; b = 8'd169;  #10 
a = 8'd15; b = 8'd170;  #10 
a = 8'd15; b = 8'd171;  #10 
a = 8'd15; b = 8'd172;  #10 
a = 8'd15; b = 8'd173;  #10 
a = 8'd15; b = 8'd174;  #10 
a = 8'd15; b = 8'd175;  #10 
a = 8'd15; b = 8'd176;  #10 
a = 8'd15; b = 8'd177;  #10 
a = 8'd15; b = 8'd178;  #10 
a = 8'd15; b = 8'd179;  #10 
a = 8'd15; b = 8'd180;  #10 
a = 8'd15; b = 8'd181;  #10 
a = 8'd15; b = 8'd182;  #10 
a = 8'd15; b = 8'd183;  #10 
a = 8'd15; b = 8'd184;  #10 
a = 8'd15; b = 8'd185;  #10 
a = 8'd15; b = 8'd186;  #10 
a = 8'd15; b = 8'd187;  #10 
a = 8'd15; b = 8'd188;  #10 
a = 8'd15; b = 8'd189;  #10 
a = 8'd15; b = 8'd190;  #10 
a = 8'd15; b = 8'd191;  #10 
a = 8'd15; b = 8'd192;  #10 
a = 8'd15; b = 8'd193;  #10 
a = 8'd15; b = 8'd194;  #10 
a = 8'd15; b = 8'd195;  #10 
a = 8'd15; b = 8'd196;  #10 
a = 8'd15; b = 8'd197;  #10 
a = 8'd15; b = 8'd198;  #10 
a = 8'd15; b = 8'd199;  #10 
a = 8'd15; b = 8'd200;  #10 
a = 8'd15; b = 8'd201;  #10 
a = 8'd15; b = 8'd202;  #10 
a = 8'd15; b = 8'd203;  #10 
a = 8'd15; b = 8'd204;  #10 
a = 8'd15; b = 8'd205;  #10 
a = 8'd15; b = 8'd206;  #10 
a = 8'd15; b = 8'd207;  #10 
a = 8'd15; b = 8'd208;  #10 
a = 8'd15; b = 8'd209;  #10 
a = 8'd15; b = 8'd210;  #10 
a = 8'd15; b = 8'd211;  #10 
a = 8'd15; b = 8'd212;  #10 
a = 8'd15; b = 8'd213;  #10 
a = 8'd15; b = 8'd214;  #10 
a = 8'd15; b = 8'd215;  #10 
a = 8'd15; b = 8'd216;  #10 
a = 8'd15; b = 8'd217;  #10 
a = 8'd15; b = 8'd218;  #10 
a = 8'd15; b = 8'd219;  #10 
a = 8'd15; b = 8'd220;  #10 
a = 8'd15; b = 8'd221;  #10 
a = 8'd15; b = 8'd222;  #10 
a = 8'd15; b = 8'd223;  #10 
a = 8'd15; b = 8'd224;  #10 
a = 8'd15; b = 8'd225;  #10 
a = 8'd15; b = 8'd226;  #10 
a = 8'd15; b = 8'd227;  #10 
a = 8'd15; b = 8'd228;  #10 
a = 8'd15; b = 8'd229;  #10 
a = 8'd15; b = 8'd230;  #10 
a = 8'd15; b = 8'd231;  #10 
a = 8'd15; b = 8'd232;  #10 
a = 8'd15; b = 8'd233;  #10 
a = 8'd15; b = 8'd234;  #10 
a = 8'd15; b = 8'd235;  #10 
a = 8'd15; b = 8'd236;  #10 
a = 8'd15; b = 8'd237;  #10 
a = 8'd15; b = 8'd238;  #10 
a = 8'd15; b = 8'd239;  #10 
a = 8'd15; b = 8'd240;  #10 
a = 8'd15; b = 8'd241;  #10 
a = 8'd15; b = 8'd242;  #10 
a = 8'd15; b = 8'd243;  #10 
a = 8'd15; b = 8'd244;  #10 
a = 8'd15; b = 8'd245;  #10 
a = 8'd15; b = 8'd246;  #10 
a = 8'd15; b = 8'd247;  #10 
a = 8'd15; b = 8'd248;  #10 
a = 8'd15; b = 8'd249;  #10 
a = 8'd15; b = 8'd250;  #10 
a = 8'd15; b = 8'd251;  #10 
a = 8'd15; b = 8'd252;  #10 
a = 8'd15; b = 8'd253;  #10 
a = 8'd15; b = 8'd254;  #10 
a = 8'd15; b = 8'd255;  #10 
a = 8'd16; b = 8'd0;  #10 
a = 8'd16; b = 8'd1;  #10 
a = 8'd16; b = 8'd2;  #10 
a = 8'd16; b = 8'd3;  #10 
a = 8'd16; b = 8'd4;  #10 
a = 8'd16; b = 8'd5;  #10 
a = 8'd16; b = 8'd6;  #10 
a = 8'd16; b = 8'd7;  #10 
a = 8'd16; b = 8'd8;  #10 
a = 8'd16; b = 8'd9;  #10 
a = 8'd16; b = 8'd10;  #10 
a = 8'd16; b = 8'd11;  #10 
a = 8'd16; b = 8'd12;  #10 
a = 8'd16; b = 8'd13;  #10 
a = 8'd16; b = 8'd14;  #10 
a = 8'd16; b = 8'd15;  #10 
a = 8'd16; b = 8'd16;  #10 
a = 8'd16; b = 8'd17;  #10 
a = 8'd16; b = 8'd18;  #10 
a = 8'd16; b = 8'd19;  #10 
a = 8'd16; b = 8'd20;  #10 
a = 8'd16; b = 8'd21;  #10 
a = 8'd16; b = 8'd22;  #10 
a = 8'd16; b = 8'd23;  #10 
a = 8'd16; b = 8'd24;  #10 
a = 8'd16; b = 8'd25;  #10 
a = 8'd16; b = 8'd26;  #10 
a = 8'd16; b = 8'd27;  #10 
a = 8'd16; b = 8'd28;  #10 
a = 8'd16; b = 8'd29;  #10 
a = 8'd16; b = 8'd30;  #10 
a = 8'd16; b = 8'd31;  #10 
a = 8'd16; b = 8'd32;  #10 
a = 8'd16; b = 8'd33;  #10 
a = 8'd16; b = 8'd34;  #10 
a = 8'd16; b = 8'd35;  #10 
a = 8'd16; b = 8'd36;  #10 
a = 8'd16; b = 8'd37;  #10 
a = 8'd16; b = 8'd38;  #10 
a = 8'd16; b = 8'd39;  #10 
a = 8'd16; b = 8'd40;  #10 
a = 8'd16; b = 8'd41;  #10 
a = 8'd16; b = 8'd42;  #10 
a = 8'd16; b = 8'd43;  #10 
a = 8'd16; b = 8'd44;  #10 
a = 8'd16; b = 8'd45;  #10 
a = 8'd16; b = 8'd46;  #10 
a = 8'd16; b = 8'd47;  #10 
a = 8'd16; b = 8'd48;  #10 
a = 8'd16; b = 8'd49;  #10 
a = 8'd16; b = 8'd50;  #10 
a = 8'd16; b = 8'd51;  #10 
a = 8'd16; b = 8'd52;  #10 
a = 8'd16; b = 8'd53;  #10 
a = 8'd16; b = 8'd54;  #10 
a = 8'd16; b = 8'd55;  #10 
a = 8'd16; b = 8'd56;  #10 
a = 8'd16; b = 8'd57;  #10 
a = 8'd16; b = 8'd58;  #10 
a = 8'd16; b = 8'd59;  #10 
a = 8'd16; b = 8'd60;  #10 
a = 8'd16; b = 8'd61;  #10 
a = 8'd16; b = 8'd62;  #10 
a = 8'd16; b = 8'd63;  #10 
a = 8'd16; b = 8'd64;  #10 
a = 8'd16; b = 8'd65;  #10 
a = 8'd16; b = 8'd66;  #10 
a = 8'd16; b = 8'd67;  #10 
a = 8'd16; b = 8'd68;  #10 
a = 8'd16; b = 8'd69;  #10 
a = 8'd16; b = 8'd70;  #10 
a = 8'd16; b = 8'd71;  #10 
a = 8'd16; b = 8'd72;  #10 
a = 8'd16; b = 8'd73;  #10 
a = 8'd16; b = 8'd74;  #10 
a = 8'd16; b = 8'd75;  #10 
a = 8'd16; b = 8'd76;  #10 
a = 8'd16; b = 8'd77;  #10 
a = 8'd16; b = 8'd78;  #10 
a = 8'd16; b = 8'd79;  #10 
a = 8'd16; b = 8'd80;  #10 
a = 8'd16; b = 8'd81;  #10 
a = 8'd16; b = 8'd82;  #10 
a = 8'd16; b = 8'd83;  #10 
a = 8'd16; b = 8'd84;  #10 
a = 8'd16; b = 8'd85;  #10 
a = 8'd16; b = 8'd86;  #10 
a = 8'd16; b = 8'd87;  #10 
a = 8'd16; b = 8'd88;  #10 
a = 8'd16; b = 8'd89;  #10 
a = 8'd16; b = 8'd90;  #10 
a = 8'd16; b = 8'd91;  #10 
a = 8'd16; b = 8'd92;  #10 
a = 8'd16; b = 8'd93;  #10 
a = 8'd16; b = 8'd94;  #10 
a = 8'd16; b = 8'd95;  #10 
a = 8'd16; b = 8'd96;  #10 
a = 8'd16; b = 8'd97;  #10 
a = 8'd16; b = 8'd98;  #10 
a = 8'd16; b = 8'd99;  #10 
a = 8'd16; b = 8'd100;  #10 
a = 8'd16; b = 8'd101;  #10 
a = 8'd16; b = 8'd102;  #10 
a = 8'd16; b = 8'd103;  #10 
a = 8'd16; b = 8'd104;  #10 
a = 8'd16; b = 8'd105;  #10 
a = 8'd16; b = 8'd106;  #10 
a = 8'd16; b = 8'd107;  #10 
a = 8'd16; b = 8'd108;  #10 
a = 8'd16; b = 8'd109;  #10 
a = 8'd16; b = 8'd110;  #10 
a = 8'd16; b = 8'd111;  #10 
a = 8'd16; b = 8'd112;  #10 
a = 8'd16; b = 8'd113;  #10 
a = 8'd16; b = 8'd114;  #10 
a = 8'd16; b = 8'd115;  #10 
a = 8'd16; b = 8'd116;  #10 
a = 8'd16; b = 8'd117;  #10 
a = 8'd16; b = 8'd118;  #10 
a = 8'd16; b = 8'd119;  #10 
a = 8'd16; b = 8'd120;  #10 
a = 8'd16; b = 8'd121;  #10 
a = 8'd16; b = 8'd122;  #10 
a = 8'd16; b = 8'd123;  #10 
a = 8'd16; b = 8'd124;  #10 
a = 8'd16; b = 8'd125;  #10 
a = 8'd16; b = 8'd126;  #10 
a = 8'd16; b = 8'd127;  #10 
a = 8'd16; b = 8'd128;  #10 
a = 8'd16; b = 8'd129;  #10 
a = 8'd16; b = 8'd130;  #10 
a = 8'd16; b = 8'd131;  #10 
a = 8'd16; b = 8'd132;  #10 
a = 8'd16; b = 8'd133;  #10 
a = 8'd16; b = 8'd134;  #10 
a = 8'd16; b = 8'd135;  #10 
a = 8'd16; b = 8'd136;  #10 
a = 8'd16; b = 8'd137;  #10 
a = 8'd16; b = 8'd138;  #10 
a = 8'd16; b = 8'd139;  #10 
a = 8'd16; b = 8'd140;  #10 
a = 8'd16; b = 8'd141;  #10 
a = 8'd16; b = 8'd142;  #10 
a = 8'd16; b = 8'd143;  #10 
a = 8'd16; b = 8'd144;  #10 
a = 8'd16; b = 8'd145;  #10 
a = 8'd16; b = 8'd146;  #10 
a = 8'd16; b = 8'd147;  #10 
a = 8'd16; b = 8'd148;  #10 
a = 8'd16; b = 8'd149;  #10 
a = 8'd16; b = 8'd150;  #10 
a = 8'd16; b = 8'd151;  #10 
a = 8'd16; b = 8'd152;  #10 
a = 8'd16; b = 8'd153;  #10 
a = 8'd16; b = 8'd154;  #10 
a = 8'd16; b = 8'd155;  #10 
a = 8'd16; b = 8'd156;  #10 
a = 8'd16; b = 8'd157;  #10 
a = 8'd16; b = 8'd158;  #10 
a = 8'd16; b = 8'd159;  #10 
a = 8'd16; b = 8'd160;  #10 
a = 8'd16; b = 8'd161;  #10 
a = 8'd16; b = 8'd162;  #10 
a = 8'd16; b = 8'd163;  #10 
a = 8'd16; b = 8'd164;  #10 
a = 8'd16; b = 8'd165;  #10 
a = 8'd16; b = 8'd166;  #10 
a = 8'd16; b = 8'd167;  #10 
a = 8'd16; b = 8'd168;  #10 
a = 8'd16; b = 8'd169;  #10 
a = 8'd16; b = 8'd170;  #10 
a = 8'd16; b = 8'd171;  #10 
a = 8'd16; b = 8'd172;  #10 
a = 8'd16; b = 8'd173;  #10 
a = 8'd16; b = 8'd174;  #10 
a = 8'd16; b = 8'd175;  #10 
a = 8'd16; b = 8'd176;  #10 
a = 8'd16; b = 8'd177;  #10 
a = 8'd16; b = 8'd178;  #10 
a = 8'd16; b = 8'd179;  #10 
a = 8'd16; b = 8'd180;  #10 
a = 8'd16; b = 8'd181;  #10 
a = 8'd16; b = 8'd182;  #10 
a = 8'd16; b = 8'd183;  #10 
a = 8'd16; b = 8'd184;  #10 
a = 8'd16; b = 8'd185;  #10 
a = 8'd16; b = 8'd186;  #10 
a = 8'd16; b = 8'd187;  #10 
a = 8'd16; b = 8'd188;  #10 
a = 8'd16; b = 8'd189;  #10 
a = 8'd16; b = 8'd190;  #10 
a = 8'd16; b = 8'd191;  #10 
a = 8'd16; b = 8'd192;  #10 
a = 8'd16; b = 8'd193;  #10 
a = 8'd16; b = 8'd194;  #10 
a = 8'd16; b = 8'd195;  #10 
a = 8'd16; b = 8'd196;  #10 
a = 8'd16; b = 8'd197;  #10 
a = 8'd16; b = 8'd198;  #10 
a = 8'd16; b = 8'd199;  #10 
a = 8'd16; b = 8'd200;  #10 
a = 8'd16; b = 8'd201;  #10 
a = 8'd16; b = 8'd202;  #10 
a = 8'd16; b = 8'd203;  #10 
a = 8'd16; b = 8'd204;  #10 
a = 8'd16; b = 8'd205;  #10 
a = 8'd16; b = 8'd206;  #10 
a = 8'd16; b = 8'd207;  #10 
a = 8'd16; b = 8'd208;  #10 
a = 8'd16; b = 8'd209;  #10 
a = 8'd16; b = 8'd210;  #10 
a = 8'd16; b = 8'd211;  #10 
a = 8'd16; b = 8'd212;  #10 
a = 8'd16; b = 8'd213;  #10 
a = 8'd16; b = 8'd214;  #10 
a = 8'd16; b = 8'd215;  #10 
a = 8'd16; b = 8'd216;  #10 
a = 8'd16; b = 8'd217;  #10 
a = 8'd16; b = 8'd218;  #10 
a = 8'd16; b = 8'd219;  #10 
a = 8'd16; b = 8'd220;  #10 
a = 8'd16; b = 8'd221;  #10 
a = 8'd16; b = 8'd222;  #10 
a = 8'd16; b = 8'd223;  #10 
a = 8'd16; b = 8'd224;  #10 
a = 8'd16; b = 8'd225;  #10 
a = 8'd16; b = 8'd226;  #10 
a = 8'd16; b = 8'd227;  #10 
a = 8'd16; b = 8'd228;  #10 
a = 8'd16; b = 8'd229;  #10 
a = 8'd16; b = 8'd230;  #10 
a = 8'd16; b = 8'd231;  #10 
a = 8'd16; b = 8'd232;  #10 
a = 8'd16; b = 8'd233;  #10 
a = 8'd16; b = 8'd234;  #10 
a = 8'd16; b = 8'd235;  #10 
a = 8'd16; b = 8'd236;  #10 
a = 8'd16; b = 8'd237;  #10 
a = 8'd16; b = 8'd238;  #10 
a = 8'd16; b = 8'd239;  #10 
a = 8'd16; b = 8'd240;  #10 
a = 8'd16; b = 8'd241;  #10 
a = 8'd16; b = 8'd242;  #10 
a = 8'd16; b = 8'd243;  #10 
a = 8'd16; b = 8'd244;  #10 
a = 8'd16; b = 8'd245;  #10 
a = 8'd16; b = 8'd246;  #10 
a = 8'd16; b = 8'd247;  #10 
a = 8'd16; b = 8'd248;  #10 
a = 8'd16; b = 8'd249;  #10 
a = 8'd16; b = 8'd250;  #10 
a = 8'd16; b = 8'd251;  #10 
a = 8'd16; b = 8'd252;  #10 
a = 8'd16; b = 8'd253;  #10 
a = 8'd16; b = 8'd254;  #10 
a = 8'd16; b = 8'd255;  #10 
a = 8'd17; b = 8'd0;  #10 
a = 8'd17; b = 8'd1;  #10 
a = 8'd17; b = 8'd2;  #10 
a = 8'd17; b = 8'd3;  #10 
a = 8'd17; b = 8'd4;  #10 
a = 8'd17; b = 8'd5;  #10 
a = 8'd17; b = 8'd6;  #10 
a = 8'd17; b = 8'd7;  #10 
a = 8'd17; b = 8'd8;  #10 
a = 8'd17; b = 8'd9;  #10 
a = 8'd17; b = 8'd10;  #10 
a = 8'd17; b = 8'd11;  #10 
a = 8'd17; b = 8'd12;  #10 
a = 8'd17; b = 8'd13;  #10 
a = 8'd17; b = 8'd14;  #10 
a = 8'd17; b = 8'd15;  #10 
a = 8'd17; b = 8'd16;  #10 
a = 8'd17; b = 8'd17;  #10 
a = 8'd17; b = 8'd18;  #10 
a = 8'd17; b = 8'd19;  #10 
a = 8'd17; b = 8'd20;  #10 
a = 8'd17; b = 8'd21;  #10 
a = 8'd17; b = 8'd22;  #10 
a = 8'd17; b = 8'd23;  #10 
a = 8'd17; b = 8'd24;  #10 
a = 8'd17; b = 8'd25;  #10 
a = 8'd17; b = 8'd26;  #10 
a = 8'd17; b = 8'd27;  #10 
a = 8'd17; b = 8'd28;  #10 
a = 8'd17; b = 8'd29;  #10 
a = 8'd17; b = 8'd30;  #10 
a = 8'd17; b = 8'd31;  #10 
a = 8'd17; b = 8'd32;  #10 
a = 8'd17; b = 8'd33;  #10 
a = 8'd17; b = 8'd34;  #10 
a = 8'd17; b = 8'd35;  #10 
a = 8'd17; b = 8'd36;  #10 
a = 8'd17; b = 8'd37;  #10 
a = 8'd17; b = 8'd38;  #10 
a = 8'd17; b = 8'd39;  #10 
a = 8'd17; b = 8'd40;  #10 
a = 8'd17; b = 8'd41;  #10 
a = 8'd17; b = 8'd42;  #10 
a = 8'd17; b = 8'd43;  #10 
a = 8'd17; b = 8'd44;  #10 
a = 8'd17; b = 8'd45;  #10 
a = 8'd17; b = 8'd46;  #10 
a = 8'd17; b = 8'd47;  #10 
a = 8'd17; b = 8'd48;  #10 
a = 8'd17; b = 8'd49;  #10 
a = 8'd17; b = 8'd50;  #10 
a = 8'd17; b = 8'd51;  #10 
a = 8'd17; b = 8'd52;  #10 
a = 8'd17; b = 8'd53;  #10 
a = 8'd17; b = 8'd54;  #10 
a = 8'd17; b = 8'd55;  #10 
a = 8'd17; b = 8'd56;  #10 
a = 8'd17; b = 8'd57;  #10 
a = 8'd17; b = 8'd58;  #10 
a = 8'd17; b = 8'd59;  #10 
a = 8'd17; b = 8'd60;  #10 
a = 8'd17; b = 8'd61;  #10 
a = 8'd17; b = 8'd62;  #10 
a = 8'd17; b = 8'd63;  #10 
a = 8'd17; b = 8'd64;  #10 
a = 8'd17; b = 8'd65;  #10 
a = 8'd17; b = 8'd66;  #10 
a = 8'd17; b = 8'd67;  #10 
a = 8'd17; b = 8'd68;  #10 
a = 8'd17; b = 8'd69;  #10 
a = 8'd17; b = 8'd70;  #10 
a = 8'd17; b = 8'd71;  #10 
a = 8'd17; b = 8'd72;  #10 
a = 8'd17; b = 8'd73;  #10 
a = 8'd17; b = 8'd74;  #10 
a = 8'd17; b = 8'd75;  #10 
a = 8'd17; b = 8'd76;  #10 
a = 8'd17; b = 8'd77;  #10 
a = 8'd17; b = 8'd78;  #10 
a = 8'd17; b = 8'd79;  #10 
a = 8'd17; b = 8'd80;  #10 
a = 8'd17; b = 8'd81;  #10 
a = 8'd17; b = 8'd82;  #10 
a = 8'd17; b = 8'd83;  #10 
a = 8'd17; b = 8'd84;  #10 
a = 8'd17; b = 8'd85;  #10 
a = 8'd17; b = 8'd86;  #10 
a = 8'd17; b = 8'd87;  #10 
a = 8'd17; b = 8'd88;  #10 
a = 8'd17; b = 8'd89;  #10 
a = 8'd17; b = 8'd90;  #10 
a = 8'd17; b = 8'd91;  #10 
a = 8'd17; b = 8'd92;  #10 
a = 8'd17; b = 8'd93;  #10 
a = 8'd17; b = 8'd94;  #10 
a = 8'd17; b = 8'd95;  #10 
a = 8'd17; b = 8'd96;  #10 
a = 8'd17; b = 8'd97;  #10 
a = 8'd17; b = 8'd98;  #10 
a = 8'd17; b = 8'd99;  #10 
a = 8'd17; b = 8'd100;  #10 
a = 8'd17; b = 8'd101;  #10 
a = 8'd17; b = 8'd102;  #10 
a = 8'd17; b = 8'd103;  #10 
a = 8'd17; b = 8'd104;  #10 
a = 8'd17; b = 8'd105;  #10 
a = 8'd17; b = 8'd106;  #10 
a = 8'd17; b = 8'd107;  #10 
a = 8'd17; b = 8'd108;  #10 
a = 8'd17; b = 8'd109;  #10 
a = 8'd17; b = 8'd110;  #10 
a = 8'd17; b = 8'd111;  #10 
a = 8'd17; b = 8'd112;  #10 
a = 8'd17; b = 8'd113;  #10 
a = 8'd17; b = 8'd114;  #10 
a = 8'd17; b = 8'd115;  #10 
a = 8'd17; b = 8'd116;  #10 
a = 8'd17; b = 8'd117;  #10 
a = 8'd17; b = 8'd118;  #10 
a = 8'd17; b = 8'd119;  #10 
a = 8'd17; b = 8'd120;  #10 
a = 8'd17; b = 8'd121;  #10 
a = 8'd17; b = 8'd122;  #10 
a = 8'd17; b = 8'd123;  #10 
a = 8'd17; b = 8'd124;  #10 
a = 8'd17; b = 8'd125;  #10 
a = 8'd17; b = 8'd126;  #10 
a = 8'd17; b = 8'd127;  #10 
a = 8'd17; b = 8'd128;  #10 
a = 8'd17; b = 8'd129;  #10 
a = 8'd17; b = 8'd130;  #10 
a = 8'd17; b = 8'd131;  #10 
a = 8'd17; b = 8'd132;  #10 
a = 8'd17; b = 8'd133;  #10 
a = 8'd17; b = 8'd134;  #10 
a = 8'd17; b = 8'd135;  #10 
a = 8'd17; b = 8'd136;  #10 
a = 8'd17; b = 8'd137;  #10 
a = 8'd17; b = 8'd138;  #10 
a = 8'd17; b = 8'd139;  #10 
a = 8'd17; b = 8'd140;  #10 
a = 8'd17; b = 8'd141;  #10 
a = 8'd17; b = 8'd142;  #10 
a = 8'd17; b = 8'd143;  #10 
a = 8'd17; b = 8'd144;  #10 
a = 8'd17; b = 8'd145;  #10 
a = 8'd17; b = 8'd146;  #10 
a = 8'd17; b = 8'd147;  #10 
a = 8'd17; b = 8'd148;  #10 
a = 8'd17; b = 8'd149;  #10 
a = 8'd17; b = 8'd150;  #10 
a = 8'd17; b = 8'd151;  #10 
a = 8'd17; b = 8'd152;  #10 
a = 8'd17; b = 8'd153;  #10 
a = 8'd17; b = 8'd154;  #10 
a = 8'd17; b = 8'd155;  #10 
a = 8'd17; b = 8'd156;  #10 
a = 8'd17; b = 8'd157;  #10 
a = 8'd17; b = 8'd158;  #10 
a = 8'd17; b = 8'd159;  #10 
a = 8'd17; b = 8'd160;  #10 
a = 8'd17; b = 8'd161;  #10 
a = 8'd17; b = 8'd162;  #10 
a = 8'd17; b = 8'd163;  #10 
a = 8'd17; b = 8'd164;  #10 
a = 8'd17; b = 8'd165;  #10 
a = 8'd17; b = 8'd166;  #10 
a = 8'd17; b = 8'd167;  #10 
a = 8'd17; b = 8'd168;  #10 
a = 8'd17; b = 8'd169;  #10 
a = 8'd17; b = 8'd170;  #10 
a = 8'd17; b = 8'd171;  #10 
a = 8'd17; b = 8'd172;  #10 
a = 8'd17; b = 8'd173;  #10 
a = 8'd17; b = 8'd174;  #10 
a = 8'd17; b = 8'd175;  #10 
a = 8'd17; b = 8'd176;  #10 
a = 8'd17; b = 8'd177;  #10 
a = 8'd17; b = 8'd178;  #10 
a = 8'd17; b = 8'd179;  #10 
a = 8'd17; b = 8'd180;  #10 
a = 8'd17; b = 8'd181;  #10 
a = 8'd17; b = 8'd182;  #10 
a = 8'd17; b = 8'd183;  #10 
a = 8'd17; b = 8'd184;  #10 
a = 8'd17; b = 8'd185;  #10 
a = 8'd17; b = 8'd186;  #10 
a = 8'd17; b = 8'd187;  #10 
a = 8'd17; b = 8'd188;  #10 
a = 8'd17; b = 8'd189;  #10 
a = 8'd17; b = 8'd190;  #10 
a = 8'd17; b = 8'd191;  #10 
a = 8'd17; b = 8'd192;  #10 
a = 8'd17; b = 8'd193;  #10 
a = 8'd17; b = 8'd194;  #10 
a = 8'd17; b = 8'd195;  #10 
a = 8'd17; b = 8'd196;  #10 
a = 8'd17; b = 8'd197;  #10 
a = 8'd17; b = 8'd198;  #10 
a = 8'd17; b = 8'd199;  #10 
a = 8'd17; b = 8'd200;  #10 
a = 8'd17; b = 8'd201;  #10 
a = 8'd17; b = 8'd202;  #10 
a = 8'd17; b = 8'd203;  #10 
a = 8'd17; b = 8'd204;  #10 
a = 8'd17; b = 8'd205;  #10 
a = 8'd17; b = 8'd206;  #10 
a = 8'd17; b = 8'd207;  #10 
a = 8'd17; b = 8'd208;  #10 
a = 8'd17; b = 8'd209;  #10 
a = 8'd17; b = 8'd210;  #10 
a = 8'd17; b = 8'd211;  #10 
a = 8'd17; b = 8'd212;  #10 
a = 8'd17; b = 8'd213;  #10 
a = 8'd17; b = 8'd214;  #10 
a = 8'd17; b = 8'd215;  #10 
a = 8'd17; b = 8'd216;  #10 
a = 8'd17; b = 8'd217;  #10 
a = 8'd17; b = 8'd218;  #10 
a = 8'd17; b = 8'd219;  #10 
a = 8'd17; b = 8'd220;  #10 
a = 8'd17; b = 8'd221;  #10 
a = 8'd17; b = 8'd222;  #10 
a = 8'd17; b = 8'd223;  #10 
a = 8'd17; b = 8'd224;  #10 
a = 8'd17; b = 8'd225;  #10 
a = 8'd17; b = 8'd226;  #10 
a = 8'd17; b = 8'd227;  #10 
a = 8'd17; b = 8'd228;  #10 
a = 8'd17; b = 8'd229;  #10 
a = 8'd17; b = 8'd230;  #10 
a = 8'd17; b = 8'd231;  #10 
a = 8'd17; b = 8'd232;  #10 
a = 8'd17; b = 8'd233;  #10 
a = 8'd17; b = 8'd234;  #10 
a = 8'd17; b = 8'd235;  #10 
a = 8'd17; b = 8'd236;  #10 
a = 8'd17; b = 8'd237;  #10 
a = 8'd17; b = 8'd238;  #10 
a = 8'd17; b = 8'd239;  #10 
a = 8'd17; b = 8'd240;  #10 
a = 8'd17; b = 8'd241;  #10 
a = 8'd17; b = 8'd242;  #10 
a = 8'd17; b = 8'd243;  #10 
a = 8'd17; b = 8'd244;  #10 
a = 8'd17; b = 8'd245;  #10 
a = 8'd17; b = 8'd246;  #10 
a = 8'd17; b = 8'd247;  #10 
a = 8'd17; b = 8'd248;  #10 
a = 8'd17; b = 8'd249;  #10 
a = 8'd17; b = 8'd250;  #10 
a = 8'd17; b = 8'd251;  #10 
a = 8'd17; b = 8'd252;  #10 
a = 8'd17; b = 8'd253;  #10 
a = 8'd17; b = 8'd254;  #10 
a = 8'd17; b = 8'd255;  #10 
a = 8'd18; b = 8'd0;  #10 
a = 8'd18; b = 8'd1;  #10 
a = 8'd18; b = 8'd2;  #10 
a = 8'd18; b = 8'd3;  #10 
a = 8'd18; b = 8'd4;  #10 
a = 8'd18; b = 8'd5;  #10 
a = 8'd18; b = 8'd6;  #10 
a = 8'd18; b = 8'd7;  #10 
a = 8'd18; b = 8'd8;  #10 
a = 8'd18; b = 8'd9;  #10 
a = 8'd18; b = 8'd10;  #10 
a = 8'd18; b = 8'd11;  #10 
a = 8'd18; b = 8'd12;  #10 
a = 8'd18; b = 8'd13;  #10 
a = 8'd18; b = 8'd14;  #10 
a = 8'd18; b = 8'd15;  #10 
a = 8'd18; b = 8'd16;  #10 
a = 8'd18; b = 8'd17;  #10 
a = 8'd18; b = 8'd18;  #10 
a = 8'd18; b = 8'd19;  #10 
a = 8'd18; b = 8'd20;  #10 
a = 8'd18; b = 8'd21;  #10 
a = 8'd18; b = 8'd22;  #10 
a = 8'd18; b = 8'd23;  #10 
a = 8'd18; b = 8'd24;  #10 
a = 8'd18; b = 8'd25;  #10 
a = 8'd18; b = 8'd26;  #10 
a = 8'd18; b = 8'd27;  #10 
a = 8'd18; b = 8'd28;  #10 
a = 8'd18; b = 8'd29;  #10 
a = 8'd18; b = 8'd30;  #10 
a = 8'd18; b = 8'd31;  #10 
a = 8'd18; b = 8'd32;  #10 
a = 8'd18; b = 8'd33;  #10 
a = 8'd18; b = 8'd34;  #10 
a = 8'd18; b = 8'd35;  #10 
a = 8'd18; b = 8'd36;  #10 
a = 8'd18; b = 8'd37;  #10 
a = 8'd18; b = 8'd38;  #10 
a = 8'd18; b = 8'd39;  #10 
a = 8'd18; b = 8'd40;  #10 
a = 8'd18; b = 8'd41;  #10 
a = 8'd18; b = 8'd42;  #10 
a = 8'd18; b = 8'd43;  #10 
a = 8'd18; b = 8'd44;  #10 
a = 8'd18; b = 8'd45;  #10 
a = 8'd18; b = 8'd46;  #10 
a = 8'd18; b = 8'd47;  #10 
a = 8'd18; b = 8'd48;  #10 
a = 8'd18; b = 8'd49;  #10 
a = 8'd18; b = 8'd50;  #10 
a = 8'd18; b = 8'd51;  #10 
a = 8'd18; b = 8'd52;  #10 
a = 8'd18; b = 8'd53;  #10 
a = 8'd18; b = 8'd54;  #10 
a = 8'd18; b = 8'd55;  #10 
a = 8'd18; b = 8'd56;  #10 
a = 8'd18; b = 8'd57;  #10 
a = 8'd18; b = 8'd58;  #10 
a = 8'd18; b = 8'd59;  #10 
a = 8'd18; b = 8'd60;  #10 
a = 8'd18; b = 8'd61;  #10 
a = 8'd18; b = 8'd62;  #10 
a = 8'd18; b = 8'd63;  #10 
a = 8'd18; b = 8'd64;  #10 
a = 8'd18; b = 8'd65;  #10 
a = 8'd18; b = 8'd66;  #10 
a = 8'd18; b = 8'd67;  #10 
a = 8'd18; b = 8'd68;  #10 
a = 8'd18; b = 8'd69;  #10 
a = 8'd18; b = 8'd70;  #10 
a = 8'd18; b = 8'd71;  #10 
a = 8'd18; b = 8'd72;  #10 
a = 8'd18; b = 8'd73;  #10 
a = 8'd18; b = 8'd74;  #10 
a = 8'd18; b = 8'd75;  #10 
a = 8'd18; b = 8'd76;  #10 
a = 8'd18; b = 8'd77;  #10 
a = 8'd18; b = 8'd78;  #10 
a = 8'd18; b = 8'd79;  #10 
a = 8'd18; b = 8'd80;  #10 
a = 8'd18; b = 8'd81;  #10 
a = 8'd18; b = 8'd82;  #10 
a = 8'd18; b = 8'd83;  #10 
a = 8'd18; b = 8'd84;  #10 
a = 8'd18; b = 8'd85;  #10 
a = 8'd18; b = 8'd86;  #10 
a = 8'd18; b = 8'd87;  #10 
a = 8'd18; b = 8'd88;  #10 
a = 8'd18; b = 8'd89;  #10 
a = 8'd18; b = 8'd90;  #10 
a = 8'd18; b = 8'd91;  #10 
a = 8'd18; b = 8'd92;  #10 
a = 8'd18; b = 8'd93;  #10 
a = 8'd18; b = 8'd94;  #10 
a = 8'd18; b = 8'd95;  #10 
a = 8'd18; b = 8'd96;  #10 
a = 8'd18; b = 8'd97;  #10 
a = 8'd18; b = 8'd98;  #10 
a = 8'd18; b = 8'd99;  #10 
a = 8'd18; b = 8'd100;  #10 
a = 8'd18; b = 8'd101;  #10 
a = 8'd18; b = 8'd102;  #10 
a = 8'd18; b = 8'd103;  #10 
a = 8'd18; b = 8'd104;  #10 
a = 8'd18; b = 8'd105;  #10 
a = 8'd18; b = 8'd106;  #10 
a = 8'd18; b = 8'd107;  #10 
a = 8'd18; b = 8'd108;  #10 
a = 8'd18; b = 8'd109;  #10 
a = 8'd18; b = 8'd110;  #10 
a = 8'd18; b = 8'd111;  #10 
a = 8'd18; b = 8'd112;  #10 
a = 8'd18; b = 8'd113;  #10 
a = 8'd18; b = 8'd114;  #10 
a = 8'd18; b = 8'd115;  #10 
a = 8'd18; b = 8'd116;  #10 
a = 8'd18; b = 8'd117;  #10 
a = 8'd18; b = 8'd118;  #10 
a = 8'd18; b = 8'd119;  #10 
a = 8'd18; b = 8'd120;  #10 
a = 8'd18; b = 8'd121;  #10 
a = 8'd18; b = 8'd122;  #10 
a = 8'd18; b = 8'd123;  #10 
a = 8'd18; b = 8'd124;  #10 
a = 8'd18; b = 8'd125;  #10 
a = 8'd18; b = 8'd126;  #10 
a = 8'd18; b = 8'd127;  #10 
a = 8'd18; b = 8'd128;  #10 
a = 8'd18; b = 8'd129;  #10 
a = 8'd18; b = 8'd130;  #10 
a = 8'd18; b = 8'd131;  #10 
a = 8'd18; b = 8'd132;  #10 
a = 8'd18; b = 8'd133;  #10 
a = 8'd18; b = 8'd134;  #10 
a = 8'd18; b = 8'd135;  #10 
a = 8'd18; b = 8'd136;  #10 
a = 8'd18; b = 8'd137;  #10 
a = 8'd18; b = 8'd138;  #10 
a = 8'd18; b = 8'd139;  #10 
a = 8'd18; b = 8'd140;  #10 
a = 8'd18; b = 8'd141;  #10 
a = 8'd18; b = 8'd142;  #10 
a = 8'd18; b = 8'd143;  #10 
a = 8'd18; b = 8'd144;  #10 
a = 8'd18; b = 8'd145;  #10 
a = 8'd18; b = 8'd146;  #10 
a = 8'd18; b = 8'd147;  #10 
a = 8'd18; b = 8'd148;  #10 
a = 8'd18; b = 8'd149;  #10 
a = 8'd18; b = 8'd150;  #10 
a = 8'd18; b = 8'd151;  #10 
a = 8'd18; b = 8'd152;  #10 
a = 8'd18; b = 8'd153;  #10 
a = 8'd18; b = 8'd154;  #10 
a = 8'd18; b = 8'd155;  #10 
a = 8'd18; b = 8'd156;  #10 
a = 8'd18; b = 8'd157;  #10 
a = 8'd18; b = 8'd158;  #10 
a = 8'd18; b = 8'd159;  #10 
a = 8'd18; b = 8'd160;  #10 
a = 8'd18; b = 8'd161;  #10 
a = 8'd18; b = 8'd162;  #10 
a = 8'd18; b = 8'd163;  #10 
a = 8'd18; b = 8'd164;  #10 
a = 8'd18; b = 8'd165;  #10 
a = 8'd18; b = 8'd166;  #10 
a = 8'd18; b = 8'd167;  #10 
a = 8'd18; b = 8'd168;  #10 
a = 8'd18; b = 8'd169;  #10 
a = 8'd18; b = 8'd170;  #10 
a = 8'd18; b = 8'd171;  #10 
a = 8'd18; b = 8'd172;  #10 
a = 8'd18; b = 8'd173;  #10 
a = 8'd18; b = 8'd174;  #10 
a = 8'd18; b = 8'd175;  #10 
a = 8'd18; b = 8'd176;  #10 
a = 8'd18; b = 8'd177;  #10 
a = 8'd18; b = 8'd178;  #10 
a = 8'd18; b = 8'd179;  #10 
a = 8'd18; b = 8'd180;  #10 
a = 8'd18; b = 8'd181;  #10 
a = 8'd18; b = 8'd182;  #10 
a = 8'd18; b = 8'd183;  #10 
a = 8'd18; b = 8'd184;  #10 
a = 8'd18; b = 8'd185;  #10 
a = 8'd18; b = 8'd186;  #10 
a = 8'd18; b = 8'd187;  #10 
a = 8'd18; b = 8'd188;  #10 
a = 8'd18; b = 8'd189;  #10 
a = 8'd18; b = 8'd190;  #10 
a = 8'd18; b = 8'd191;  #10 
a = 8'd18; b = 8'd192;  #10 
a = 8'd18; b = 8'd193;  #10 
a = 8'd18; b = 8'd194;  #10 
a = 8'd18; b = 8'd195;  #10 
a = 8'd18; b = 8'd196;  #10 
a = 8'd18; b = 8'd197;  #10 
a = 8'd18; b = 8'd198;  #10 
a = 8'd18; b = 8'd199;  #10 
a = 8'd18; b = 8'd200;  #10 
a = 8'd18; b = 8'd201;  #10 
a = 8'd18; b = 8'd202;  #10 
a = 8'd18; b = 8'd203;  #10 
a = 8'd18; b = 8'd204;  #10 
a = 8'd18; b = 8'd205;  #10 
a = 8'd18; b = 8'd206;  #10 
a = 8'd18; b = 8'd207;  #10 
a = 8'd18; b = 8'd208;  #10 
a = 8'd18; b = 8'd209;  #10 
a = 8'd18; b = 8'd210;  #10 
a = 8'd18; b = 8'd211;  #10 
a = 8'd18; b = 8'd212;  #10 
a = 8'd18; b = 8'd213;  #10 
a = 8'd18; b = 8'd214;  #10 
a = 8'd18; b = 8'd215;  #10 
a = 8'd18; b = 8'd216;  #10 
a = 8'd18; b = 8'd217;  #10 
a = 8'd18; b = 8'd218;  #10 
a = 8'd18; b = 8'd219;  #10 
a = 8'd18; b = 8'd220;  #10 
a = 8'd18; b = 8'd221;  #10 
a = 8'd18; b = 8'd222;  #10 
a = 8'd18; b = 8'd223;  #10 
a = 8'd18; b = 8'd224;  #10 
a = 8'd18; b = 8'd225;  #10 
a = 8'd18; b = 8'd226;  #10 
a = 8'd18; b = 8'd227;  #10 
a = 8'd18; b = 8'd228;  #10 
a = 8'd18; b = 8'd229;  #10 
a = 8'd18; b = 8'd230;  #10 
a = 8'd18; b = 8'd231;  #10 
a = 8'd18; b = 8'd232;  #10 
a = 8'd18; b = 8'd233;  #10 
a = 8'd18; b = 8'd234;  #10 
a = 8'd18; b = 8'd235;  #10 
a = 8'd18; b = 8'd236;  #10 
a = 8'd18; b = 8'd237;  #10 
a = 8'd18; b = 8'd238;  #10 
a = 8'd18; b = 8'd239;  #10 
a = 8'd18; b = 8'd240;  #10 
a = 8'd18; b = 8'd241;  #10 
a = 8'd18; b = 8'd242;  #10 
a = 8'd18; b = 8'd243;  #10 
a = 8'd18; b = 8'd244;  #10 
a = 8'd18; b = 8'd245;  #10 
a = 8'd18; b = 8'd246;  #10 
a = 8'd18; b = 8'd247;  #10 
a = 8'd18; b = 8'd248;  #10 
a = 8'd18; b = 8'd249;  #10 
a = 8'd18; b = 8'd250;  #10 
a = 8'd18; b = 8'd251;  #10 
a = 8'd18; b = 8'd252;  #10 
a = 8'd18; b = 8'd253;  #10 
a = 8'd18; b = 8'd254;  #10 
a = 8'd18; b = 8'd255;  #10 
a = 8'd19; b = 8'd0;  #10 
a = 8'd19; b = 8'd1;  #10 
a = 8'd19; b = 8'd2;  #10 
a = 8'd19; b = 8'd3;  #10 
a = 8'd19; b = 8'd4;  #10 
a = 8'd19; b = 8'd5;  #10 
a = 8'd19; b = 8'd6;  #10 
a = 8'd19; b = 8'd7;  #10 
a = 8'd19; b = 8'd8;  #10 
a = 8'd19; b = 8'd9;  #10 
a = 8'd19; b = 8'd10;  #10 
a = 8'd19; b = 8'd11;  #10 
a = 8'd19; b = 8'd12;  #10 
a = 8'd19; b = 8'd13;  #10 
a = 8'd19; b = 8'd14;  #10 
a = 8'd19; b = 8'd15;  #10 
a = 8'd19; b = 8'd16;  #10 
a = 8'd19; b = 8'd17;  #10 
a = 8'd19; b = 8'd18;  #10 
a = 8'd19; b = 8'd19;  #10 
a = 8'd19; b = 8'd20;  #10 
a = 8'd19; b = 8'd21;  #10 
a = 8'd19; b = 8'd22;  #10 
a = 8'd19; b = 8'd23;  #10 
a = 8'd19; b = 8'd24;  #10 
a = 8'd19; b = 8'd25;  #10 
a = 8'd19; b = 8'd26;  #10 
a = 8'd19; b = 8'd27;  #10 
a = 8'd19; b = 8'd28;  #10 
a = 8'd19; b = 8'd29;  #10 
a = 8'd19; b = 8'd30;  #10 
a = 8'd19; b = 8'd31;  #10 
a = 8'd19; b = 8'd32;  #10 
a = 8'd19; b = 8'd33;  #10 
a = 8'd19; b = 8'd34;  #10 
a = 8'd19; b = 8'd35;  #10 
a = 8'd19; b = 8'd36;  #10 
a = 8'd19; b = 8'd37;  #10 
a = 8'd19; b = 8'd38;  #10 
a = 8'd19; b = 8'd39;  #10 
a = 8'd19; b = 8'd40;  #10 
a = 8'd19; b = 8'd41;  #10 
a = 8'd19; b = 8'd42;  #10 
a = 8'd19; b = 8'd43;  #10 
a = 8'd19; b = 8'd44;  #10 
a = 8'd19; b = 8'd45;  #10 
a = 8'd19; b = 8'd46;  #10 
a = 8'd19; b = 8'd47;  #10 
a = 8'd19; b = 8'd48;  #10 
a = 8'd19; b = 8'd49;  #10 
a = 8'd19; b = 8'd50;  #10 
a = 8'd19; b = 8'd51;  #10 
a = 8'd19; b = 8'd52;  #10 
a = 8'd19; b = 8'd53;  #10 
a = 8'd19; b = 8'd54;  #10 
a = 8'd19; b = 8'd55;  #10 
a = 8'd19; b = 8'd56;  #10 
a = 8'd19; b = 8'd57;  #10 
a = 8'd19; b = 8'd58;  #10 
a = 8'd19; b = 8'd59;  #10 
a = 8'd19; b = 8'd60;  #10 
a = 8'd19; b = 8'd61;  #10 
a = 8'd19; b = 8'd62;  #10 
a = 8'd19; b = 8'd63;  #10 
a = 8'd19; b = 8'd64;  #10 
a = 8'd19; b = 8'd65;  #10 
a = 8'd19; b = 8'd66;  #10 
a = 8'd19; b = 8'd67;  #10 
a = 8'd19; b = 8'd68;  #10 
a = 8'd19; b = 8'd69;  #10 
a = 8'd19; b = 8'd70;  #10 
a = 8'd19; b = 8'd71;  #10 
a = 8'd19; b = 8'd72;  #10 
a = 8'd19; b = 8'd73;  #10 
a = 8'd19; b = 8'd74;  #10 
a = 8'd19; b = 8'd75;  #10 
a = 8'd19; b = 8'd76;  #10 
a = 8'd19; b = 8'd77;  #10 
a = 8'd19; b = 8'd78;  #10 
a = 8'd19; b = 8'd79;  #10 
a = 8'd19; b = 8'd80;  #10 
a = 8'd19; b = 8'd81;  #10 
a = 8'd19; b = 8'd82;  #10 
a = 8'd19; b = 8'd83;  #10 
a = 8'd19; b = 8'd84;  #10 
a = 8'd19; b = 8'd85;  #10 
a = 8'd19; b = 8'd86;  #10 
a = 8'd19; b = 8'd87;  #10 
a = 8'd19; b = 8'd88;  #10 
a = 8'd19; b = 8'd89;  #10 
a = 8'd19; b = 8'd90;  #10 
a = 8'd19; b = 8'd91;  #10 
a = 8'd19; b = 8'd92;  #10 
a = 8'd19; b = 8'd93;  #10 
a = 8'd19; b = 8'd94;  #10 
a = 8'd19; b = 8'd95;  #10 
a = 8'd19; b = 8'd96;  #10 
a = 8'd19; b = 8'd97;  #10 
a = 8'd19; b = 8'd98;  #10 
a = 8'd19; b = 8'd99;  #10 
a = 8'd19; b = 8'd100;  #10 
a = 8'd19; b = 8'd101;  #10 
a = 8'd19; b = 8'd102;  #10 
a = 8'd19; b = 8'd103;  #10 
a = 8'd19; b = 8'd104;  #10 
a = 8'd19; b = 8'd105;  #10 
a = 8'd19; b = 8'd106;  #10 
a = 8'd19; b = 8'd107;  #10 
a = 8'd19; b = 8'd108;  #10 
a = 8'd19; b = 8'd109;  #10 
a = 8'd19; b = 8'd110;  #10 
a = 8'd19; b = 8'd111;  #10 
a = 8'd19; b = 8'd112;  #10 
a = 8'd19; b = 8'd113;  #10 
a = 8'd19; b = 8'd114;  #10 
a = 8'd19; b = 8'd115;  #10 
a = 8'd19; b = 8'd116;  #10 
a = 8'd19; b = 8'd117;  #10 
a = 8'd19; b = 8'd118;  #10 
a = 8'd19; b = 8'd119;  #10 
a = 8'd19; b = 8'd120;  #10 
a = 8'd19; b = 8'd121;  #10 
a = 8'd19; b = 8'd122;  #10 
a = 8'd19; b = 8'd123;  #10 
a = 8'd19; b = 8'd124;  #10 
a = 8'd19; b = 8'd125;  #10 
a = 8'd19; b = 8'd126;  #10 
a = 8'd19; b = 8'd127;  #10 
a = 8'd19; b = 8'd128;  #10 
a = 8'd19; b = 8'd129;  #10 
a = 8'd19; b = 8'd130;  #10 
a = 8'd19; b = 8'd131;  #10 
a = 8'd19; b = 8'd132;  #10 
a = 8'd19; b = 8'd133;  #10 
a = 8'd19; b = 8'd134;  #10 
a = 8'd19; b = 8'd135;  #10 
a = 8'd19; b = 8'd136;  #10 
a = 8'd19; b = 8'd137;  #10 
a = 8'd19; b = 8'd138;  #10 
a = 8'd19; b = 8'd139;  #10 
a = 8'd19; b = 8'd140;  #10 
a = 8'd19; b = 8'd141;  #10 
a = 8'd19; b = 8'd142;  #10 
a = 8'd19; b = 8'd143;  #10 
a = 8'd19; b = 8'd144;  #10 
a = 8'd19; b = 8'd145;  #10 
a = 8'd19; b = 8'd146;  #10 
a = 8'd19; b = 8'd147;  #10 
a = 8'd19; b = 8'd148;  #10 
a = 8'd19; b = 8'd149;  #10 
a = 8'd19; b = 8'd150;  #10 
a = 8'd19; b = 8'd151;  #10 
a = 8'd19; b = 8'd152;  #10 
a = 8'd19; b = 8'd153;  #10 
a = 8'd19; b = 8'd154;  #10 
a = 8'd19; b = 8'd155;  #10 
a = 8'd19; b = 8'd156;  #10 
a = 8'd19; b = 8'd157;  #10 
a = 8'd19; b = 8'd158;  #10 
a = 8'd19; b = 8'd159;  #10 
a = 8'd19; b = 8'd160;  #10 
a = 8'd19; b = 8'd161;  #10 
a = 8'd19; b = 8'd162;  #10 
a = 8'd19; b = 8'd163;  #10 
a = 8'd19; b = 8'd164;  #10 
a = 8'd19; b = 8'd165;  #10 
a = 8'd19; b = 8'd166;  #10 
a = 8'd19; b = 8'd167;  #10 
a = 8'd19; b = 8'd168;  #10 
a = 8'd19; b = 8'd169;  #10 
a = 8'd19; b = 8'd170;  #10 
a = 8'd19; b = 8'd171;  #10 
a = 8'd19; b = 8'd172;  #10 
a = 8'd19; b = 8'd173;  #10 
a = 8'd19; b = 8'd174;  #10 
a = 8'd19; b = 8'd175;  #10 
a = 8'd19; b = 8'd176;  #10 
a = 8'd19; b = 8'd177;  #10 
a = 8'd19; b = 8'd178;  #10 
a = 8'd19; b = 8'd179;  #10 
a = 8'd19; b = 8'd180;  #10 
a = 8'd19; b = 8'd181;  #10 
a = 8'd19; b = 8'd182;  #10 
a = 8'd19; b = 8'd183;  #10 
a = 8'd19; b = 8'd184;  #10 
a = 8'd19; b = 8'd185;  #10 
a = 8'd19; b = 8'd186;  #10 
a = 8'd19; b = 8'd187;  #10 
a = 8'd19; b = 8'd188;  #10 
a = 8'd19; b = 8'd189;  #10 
a = 8'd19; b = 8'd190;  #10 
a = 8'd19; b = 8'd191;  #10 
a = 8'd19; b = 8'd192;  #10 
a = 8'd19; b = 8'd193;  #10 
a = 8'd19; b = 8'd194;  #10 
a = 8'd19; b = 8'd195;  #10 
a = 8'd19; b = 8'd196;  #10 
a = 8'd19; b = 8'd197;  #10 
a = 8'd19; b = 8'd198;  #10 
a = 8'd19; b = 8'd199;  #10 
a = 8'd19; b = 8'd200;  #10 
a = 8'd19; b = 8'd201;  #10 
a = 8'd19; b = 8'd202;  #10 
a = 8'd19; b = 8'd203;  #10 
a = 8'd19; b = 8'd204;  #10 
a = 8'd19; b = 8'd205;  #10 
a = 8'd19; b = 8'd206;  #10 
a = 8'd19; b = 8'd207;  #10 
a = 8'd19; b = 8'd208;  #10 
a = 8'd19; b = 8'd209;  #10 
a = 8'd19; b = 8'd210;  #10 
a = 8'd19; b = 8'd211;  #10 
a = 8'd19; b = 8'd212;  #10 
a = 8'd19; b = 8'd213;  #10 
a = 8'd19; b = 8'd214;  #10 
a = 8'd19; b = 8'd215;  #10 
a = 8'd19; b = 8'd216;  #10 
a = 8'd19; b = 8'd217;  #10 
a = 8'd19; b = 8'd218;  #10 
a = 8'd19; b = 8'd219;  #10 
a = 8'd19; b = 8'd220;  #10 
a = 8'd19; b = 8'd221;  #10 
a = 8'd19; b = 8'd222;  #10 
a = 8'd19; b = 8'd223;  #10 
a = 8'd19; b = 8'd224;  #10 
a = 8'd19; b = 8'd225;  #10 
a = 8'd19; b = 8'd226;  #10 
a = 8'd19; b = 8'd227;  #10 
a = 8'd19; b = 8'd228;  #10 
a = 8'd19; b = 8'd229;  #10 
a = 8'd19; b = 8'd230;  #10 
a = 8'd19; b = 8'd231;  #10 
a = 8'd19; b = 8'd232;  #10 
a = 8'd19; b = 8'd233;  #10 
a = 8'd19; b = 8'd234;  #10 
a = 8'd19; b = 8'd235;  #10 
a = 8'd19; b = 8'd236;  #10 
a = 8'd19; b = 8'd237;  #10 
a = 8'd19; b = 8'd238;  #10 
a = 8'd19; b = 8'd239;  #10 
a = 8'd19; b = 8'd240;  #10 
a = 8'd19; b = 8'd241;  #10 
a = 8'd19; b = 8'd242;  #10 
a = 8'd19; b = 8'd243;  #10 
a = 8'd19; b = 8'd244;  #10 
a = 8'd19; b = 8'd245;  #10 
a = 8'd19; b = 8'd246;  #10 
a = 8'd19; b = 8'd247;  #10 
a = 8'd19; b = 8'd248;  #10 
a = 8'd19; b = 8'd249;  #10 
a = 8'd19; b = 8'd250;  #10 
a = 8'd19; b = 8'd251;  #10 
a = 8'd19; b = 8'd252;  #10 
a = 8'd19; b = 8'd253;  #10 
a = 8'd19; b = 8'd254;  #10 
a = 8'd19; b = 8'd255;  #10 
a = 8'd20; b = 8'd0;  #10 
a = 8'd20; b = 8'd1;  #10 
a = 8'd20; b = 8'd2;  #10 
a = 8'd20; b = 8'd3;  #10 
a = 8'd20; b = 8'd4;  #10 
a = 8'd20; b = 8'd5;  #10 
a = 8'd20; b = 8'd6;  #10 
a = 8'd20; b = 8'd7;  #10 
a = 8'd20; b = 8'd8;  #10 
a = 8'd20; b = 8'd9;  #10 
a = 8'd20; b = 8'd10;  #10 
a = 8'd20; b = 8'd11;  #10 
a = 8'd20; b = 8'd12;  #10 
a = 8'd20; b = 8'd13;  #10 
a = 8'd20; b = 8'd14;  #10 
a = 8'd20; b = 8'd15;  #10 
a = 8'd20; b = 8'd16;  #10 
a = 8'd20; b = 8'd17;  #10 
a = 8'd20; b = 8'd18;  #10 
a = 8'd20; b = 8'd19;  #10 
a = 8'd20; b = 8'd20;  #10 
a = 8'd20; b = 8'd21;  #10 
a = 8'd20; b = 8'd22;  #10 
a = 8'd20; b = 8'd23;  #10 
a = 8'd20; b = 8'd24;  #10 
a = 8'd20; b = 8'd25;  #10 
a = 8'd20; b = 8'd26;  #10 
a = 8'd20; b = 8'd27;  #10 
a = 8'd20; b = 8'd28;  #10 
a = 8'd20; b = 8'd29;  #10 
a = 8'd20; b = 8'd30;  #10 
a = 8'd20; b = 8'd31;  #10 
a = 8'd20; b = 8'd32;  #10 
a = 8'd20; b = 8'd33;  #10 
a = 8'd20; b = 8'd34;  #10 
a = 8'd20; b = 8'd35;  #10 
a = 8'd20; b = 8'd36;  #10 
a = 8'd20; b = 8'd37;  #10 
a = 8'd20; b = 8'd38;  #10 
a = 8'd20; b = 8'd39;  #10 
a = 8'd20; b = 8'd40;  #10 
a = 8'd20; b = 8'd41;  #10 
a = 8'd20; b = 8'd42;  #10 
a = 8'd20; b = 8'd43;  #10 
a = 8'd20; b = 8'd44;  #10 
a = 8'd20; b = 8'd45;  #10 
a = 8'd20; b = 8'd46;  #10 
a = 8'd20; b = 8'd47;  #10 
a = 8'd20; b = 8'd48;  #10 
a = 8'd20; b = 8'd49;  #10 
a = 8'd20; b = 8'd50;  #10 
a = 8'd20; b = 8'd51;  #10 
a = 8'd20; b = 8'd52;  #10 
a = 8'd20; b = 8'd53;  #10 
a = 8'd20; b = 8'd54;  #10 
a = 8'd20; b = 8'd55;  #10 
a = 8'd20; b = 8'd56;  #10 
a = 8'd20; b = 8'd57;  #10 
a = 8'd20; b = 8'd58;  #10 
a = 8'd20; b = 8'd59;  #10 
a = 8'd20; b = 8'd60;  #10 
a = 8'd20; b = 8'd61;  #10 
a = 8'd20; b = 8'd62;  #10 
a = 8'd20; b = 8'd63;  #10 
a = 8'd20; b = 8'd64;  #10 
a = 8'd20; b = 8'd65;  #10 
a = 8'd20; b = 8'd66;  #10 
a = 8'd20; b = 8'd67;  #10 
a = 8'd20; b = 8'd68;  #10 
a = 8'd20; b = 8'd69;  #10 
a = 8'd20; b = 8'd70;  #10 
a = 8'd20; b = 8'd71;  #10 
a = 8'd20; b = 8'd72;  #10 
a = 8'd20; b = 8'd73;  #10 
a = 8'd20; b = 8'd74;  #10 
a = 8'd20; b = 8'd75;  #10 
a = 8'd20; b = 8'd76;  #10 
a = 8'd20; b = 8'd77;  #10 
a = 8'd20; b = 8'd78;  #10 
a = 8'd20; b = 8'd79;  #10 
a = 8'd20; b = 8'd80;  #10 
a = 8'd20; b = 8'd81;  #10 
a = 8'd20; b = 8'd82;  #10 
a = 8'd20; b = 8'd83;  #10 
a = 8'd20; b = 8'd84;  #10 
a = 8'd20; b = 8'd85;  #10 
a = 8'd20; b = 8'd86;  #10 
a = 8'd20; b = 8'd87;  #10 
a = 8'd20; b = 8'd88;  #10 
a = 8'd20; b = 8'd89;  #10 
a = 8'd20; b = 8'd90;  #10 
a = 8'd20; b = 8'd91;  #10 
a = 8'd20; b = 8'd92;  #10 
a = 8'd20; b = 8'd93;  #10 
a = 8'd20; b = 8'd94;  #10 
a = 8'd20; b = 8'd95;  #10 
a = 8'd20; b = 8'd96;  #10 
a = 8'd20; b = 8'd97;  #10 
a = 8'd20; b = 8'd98;  #10 
a = 8'd20; b = 8'd99;  #10 
a = 8'd20; b = 8'd100;  #10 
a = 8'd20; b = 8'd101;  #10 
a = 8'd20; b = 8'd102;  #10 
a = 8'd20; b = 8'd103;  #10 
a = 8'd20; b = 8'd104;  #10 
a = 8'd20; b = 8'd105;  #10 
a = 8'd20; b = 8'd106;  #10 
a = 8'd20; b = 8'd107;  #10 
a = 8'd20; b = 8'd108;  #10 
a = 8'd20; b = 8'd109;  #10 
a = 8'd20; b = 8'd110;  #10 
a = 8'd20; b = 8'd111;  #10 
a = 8'd20; b = 8'd112;  #10 
a = 8'd20; b = 8'd113;  #10 
a = 8'd20; b = 8'd114;  #10 
a = 8'd20; b = 8'd115;  #10 
a = 8'd20; b = 8'd116;  #10 
a = 8'd20; b = 8'd117;  #10 
a = 8'd20; b = 8'd118;  #10 
a = 8'd20; b = 8'd119;  #10 
a = 8'd20; b = 8'd120;  #10 
a = 8'd20; b = 8'd121;  #10 
a = 8'd20; b = 8'd122;  #10 
a = 8'd20; b = 8'd123;  #10 
a = 8'd20; b = 8'd124;  #10 
a = 8'd20; b = 8'd125;  #10 
a = 8'd20; b = 8'd126;  #10 
a = 8'd20; b = 8'd127;  #10 
a = 8'd20; b = 8'd128;  #10 
a = 8'd20; b = 8'd129;  #10 
a = 8'd20; b = 8'd130;  #10 
a = 8'd20; b = 8'd131;  #10 
a = 8'd20; b = 8'd132;  #10 
a = 8'd20; b = 8'd133;  #10 
a = 8'd20; b = 8'd134;  #10 
a = 8'd20; b = 8'd135;  #10 
a = 8'd20; b = 8'd136;  #10 
a = 8'd20; b = 8'd137;  #10 
a = 8'd20; b = 8'd138;  #10 
a = 8'd20; b = 8'd139;  #10 
a = 8'd20; b = 8'd140;  #10 
a = 8'd20; b = 8'd141;  #10 
a = 8'd20; b = 8'd142;  #10 
a = 8'd20; b = 8'd143;  #10 
a = 8'd20; b = 8'd144;  #10 
a = 8'd20; b = 8'd145;  #10 
a = 8'd20; b = 8'd146;  #10 
a = 8'd20; b = 8'd147;  #10 
a = 8'd20; b = 8'd148;  #10 
a = 8'd20; b = 8'd149;  #10 
a = 8'd20; b = 8'd150;  #10 
a = 8'd20; b = 8'd151;  #10 
a = 8'd20; b = 8'd152;  #10 
a = 8'd20; b = 8'd153;  #10 
a = 8'd20; b = 8'd154;  #10 
a = 8'd20; b = 8'd155;  #10 
a = 8'd20; b = 8'd156;  #10 
a = 8'd20; b = 8'd157;  #10 
a = 8'd20; b = 8'd158;  #10 
a = 8'd20; b = 8'd159;  #10 
a = 8'd20; b = 8'd160;  #10 
a = 8'd20; b = 8'd161;  #10 
a = 8'd20; b = 8'd162;  #10 
a = 8'd20; b = 8'd163;  #10 
a = 8'd20; b = 8'd164;  #10 
a = 8'd20; b = 8'd165;  #10 
a = 8'd20; b = 8'd166;  #10 
a = 8'd20; b = 8'd167;  #10 
a = 8'd20; b = 8'd168;  #10 
a = 8'd20; b = 8'd169;  #10 
a = 8'd20; b = 8'd170;  #10 
a = 8'd20; b = 8'd171;  #10 
a = 8'd20; b = 8'd172;  #10 
a = 8'd20; b = 8'd173;  #10 
a = 8'd20; b = 8'd174;  #10 
a = 8'd20; b = 8'd175;  #10 
a = 8'd20; b = 8'd176;  #10 
a = 8'd20; b = 8'd177;  #10 
a = 8'd20; b = 8'd178;  #10 
a = 8'd20; b = 8'd179;  #10 
a = 8'd20; b = 8'd180;  #10 
a = 8'd20; b = 8'd181;  #10 
a = 8'd20; b = 8'd182;  #10 
a = 8'd20; b = 8'd183;  #10 
a = 8'd20; b = 8'd184;  #10 
a = 8'd20; b = 8'd185;  #10 
a = 8'd20; b = 8'd186;  #10 
a = 8'd20; b = 8'd187;  #10 
a = 8'd20; b = 8'd188;  #10 
a = 8'd20; b = 8'd189;  #10 
a = 8'd20; b = 8'd190;  #10 
a = 8'd20; b = 8'd191;  #10 
a = 8'd20; b = 8'd192;  #10 
a = 8'd20; b = 8'd193;  #10 
a = 8'd20; b = 8'd194;  #10 
a = 8'd20; b = 8'd195;  #10 
a = 8'd20; b = 8'd196;  #10 
a = 8'd20; b = 8'd197;  #10 
a = 8'd20; b = 8'd198;  #10 
a = 8'd20; b = 8'd199;  #10 
a = 8'd20; b = 8'd200;  #10 
a = 8'd20; b = 8'd201;  #10 
a = 8'd20; b = 8'd202;  #10 
a = 8'd20; b = 8'd203;  #10 
a = 8'd20; b = 8'd204;  #10 
a = 8'd20; b = 8'd205;  #10 
a = 8'd20; b = 8'd206;  #10 
a = 8'd20; b = 8'd207;  #10 
a = 8'd20; b = 8'd208;  #10 
a = 8'd20; b = 8'd209;  #10 
a = 8'd20; b = 8'd210;  #10 
a = 8'd20; b = 8'd211;  #10 
a = 8'd20; b = 8'd212;  #10 
a = 8'd20; b = 8'd213;  #10 
a = 8'd20; b = 8'd214;  #10 
a = 8'd20; b = 8'd215;  #10 
a = 8'd20; b = 8'd216;  #10 
a = 8'd20; b = 8'd217;  #10 
a = 8'd20; b = 8'd218;  #10 
a = 8'd20; b = 8'd219;  #10 
a = 8'd20; b = 8'd220;  #10 
a = 8'd20; b = 8'd221;  #10 
a = 8'd20; b = 8'd222;  #10 
a = 8'd20; b = 8'd223;  #10 
a = 8'd20; b = 8'd224;  #10 
a = 8'd20; b = 8'd225;  #10 
a = 8'd20; b = 8'd226;  #10 
a = 8'd20; b = 8'd227;  #10 
a = 8'd20; b = 8'd228;  #10 
a = 8'd20; b = 8'd229;  #10 
a = 8'd20; b = 8'd230;  #10 
a = 8'd20; b = 8'd231;  #10 
a = 8'd20; b = 8'd232;  #10 
a = 8'd20; b = 8'd233;  #10 
a = 8'd20; b = 8'd234;  #10 
a = 8'd20; b = 8'd235;  #10 
a = 8'd20; b = 8'd236;  #10 
a = 8'd20; b = 8'd237;  #10 
a = 8'd20; b = 8'd238;  #10 
a = 8'd20; b = 8'd239;  #10 
a = 8'd20; b = 8'd240;  #10 
a = 8'd20; b = 8'd241;  #10 
a = 8'd20; b = 8'd242;  #10 
a = 8'd20; b = 8'd243;  #10 
a = 8'd20; b = 8'd244;  #10 
a = 8'd20; b = 8'd245;  #10 
a = 8'd20; b = 8'd246;  #10 
a = 8'd20; b = 8'd247;  #10 
a = 8'd20; b = 8'd248;  #10 
a = 8'd20; b = 8'd249;  #10 
a = 8'd20; b = 8'd250;  #10 
a = 8'd20; b = 8'd251;  #10 
a = 8'd20; b = 8'd252;  #10 
a = 8'd20; b = 8'd253;  #10 
a = 8'd20; b = 8'd254;  #10 
a = 8'd20; b = 8'd255;  #10 
a = 8'd21; b = 8'd0;  #10 
a = 8'd21; b = 8'd1;  #10 
a = 8'd21; b = 8'd2;  #10 
a = 8'd21; b = 8'd3;  #10 
a = 8'd21; b = 8'd4;  #10 
a = 8'd21; b = 8'd5;  #10 
a = 8'd21; b = 8'd6;  #10 
a = 8'd21; b = 8'd7;  #10 
a = 8'd21; b = 8'd8;  #10 
a = 8'd21; b = 8'd9;  #10 
a = 8'd21; b = 8'd10;  #10 
a = 8'd21; b = 8'd11;  #10 
a = 8'd21; b = 8'd12;  #10 
a = 8'd21; b = 8'd13;  #10 
a = 8'd21; b = 8'd14;  #10 
a = 8'd21; b = 8'd15;  #10 
a = 8'd21; b = 8'd16;  #10 
a = 8'd21; b = 8'd17;  #10 
a = 8'd21; b = 8'd18;  #10 
a = 8'd21; b = 8'd19;  #10 
a = 8'd21; b = 8'd20;  #10 
a = 8'd21; b = 8'd21;  #10 
a = 8'd21; b = 8'd22;  #10 
a = 8'd21; b = 8'd23;  #10 
a = 8'd21; b = 8'd24;  #10 
a = 8'd21; b = 8'd25;  #10 
a = 8'd21; b = 8'd26;  #10 
a = 8'd21; b = 8'd27;  #10 
a = 8'd21; b = 8'd28;  #10 
a = 8'd21; b = 8'd29;  #10 
a = 8'd21; b = 8'd30;  #10 
a = 8'd21; b = 8'd31;  #10 
a = 8'd21; b = 8'd32;  #10 
a = 8'd21; b = 8'd33;  #10 
a = 8'd21; b = 8'd34;  #10 
a = 8'd21; b = 8'd35;  #10 
a = 8'd21; b = 8'd36;  #10 
a = 8'd21; b = 8'd37;  #10 
a = 8'd21; b = 8'd38;  #10 
a = 8'd21; b = 8'd39;  #10 
a = 8'd21; b = 8'd40;  #10 
a = 8'd21; b = 8'd41;  #10 
a = 8'd21; b = 8'd42;  #10 
a = 8'd21; b = 8'd43;  #10 
a = 8'd21; b = 8'd44;  #10 
a = 8'd21; b = 8'd45;  #10 
a = 8'd21; b = 8'd46;  #10 
a = 8'd21; b = 8'd47;  #10 
a = 8'd21; b = 8'd48;  #10 
a = 8'd21; b = 8'd49;  #10 
a = 8'd21; b = 8'd50;  #10 
a = 8'd21; b = 8'd51;  #10 
a = 8'd21; b = 8'd52;  #10 
a = 8'd21; b = 8'd53;  #10 
a = 8'd21; b = 8'd54;  #10 
a = 8'd21; b = 8'd55;  #10 
a = 8'd21; b = 8'd56;  #10 
a = 8'd21; b = 8'd57;  #10 
a = 8'd21; b = 8'd58;  #10 
a = 8'd21; b = 8'd59;  #10 
a = 8'd21; b = 8'd60;  #10 
a = 8'd21; b = 8'd61;  #10 
a = 8'd21; b = 8'd62;  #10 
a = 8'd21; b = 8'd63;  #10 
a = 8'd21; b = 8'd64;  #10 
a = 8'd21; b = 8'd65;  #10 
a = 8'd21; b = 8'd66;  #10 
a = 8'd21; b = 8'd67;  #10 
a = 8'd21; b = 8'd68;  #10 
a = 8'd21; b = 8'd69;  #10 
a = 8'd21; b = 8'd70;  #10 
a = 8'd21; b = 8'd71;  #10 
a = 8'd21; b = 8'd72;  #10 
a = 8'd21; b = 8'd73;  #10 
a = 8'd21; b = 8'd74;  #10 
a = 8'd21; b = 8'd75;  #10 
a = 8'd21; b = 8'd76;  #10 
a = 8'd21; b = 8'd77;  #10 
a = 8'd21; b = 8'd78;  #10 
a = 8'd21; b = 8'd79;  #10 
a = 8'd21; b = 8'd80;  #10 
a = 8'd21; b = 8'd81;  #10 
a = 8'd21; b = 8'd82;  #10 
a = 8'd21; b = 8'd83;  #10 
a = 8'd21; b = 8'd84;  #10 
a = 8'd21; b = 8'd85;  #10 
a = 8'd21; b = 8'd86;  #10 
a = 8'd21; b = 8'd87;  #10 
a = 8'd21; b = 8'd88;  #10 
a = 8'd21; b = 8'd89;  #10 
a = 8'd21; b = 8'd90;  #10 
a = 8'd21; b = 8'd91;  #10 
a = 8'd21; b = 8'd92;  #10 
a = 8'd21; b = 8'd93;  #10 
a = 8'd21; b = 8'd94;  #10 
a = 8'd21; b = 8'd95;  #10 
a = 8'd21; b = 8'd96;  #10 
a = 8'd21; b = 8'd97;  #10 
a = 8'd21; b = 8'd98;  #10 
a = 8'd21; b = 8'd99;  #10 
a = 8'd21; b = 8'd100;  #10 
a = 8'd21; b = 8'd101;  #10 
a = 8'd21; b = 8'd102;  #10 
a = 8'd21; b = 8'd103;  #10 
a = 8'd21; b = 8'd104;  #10 
a = 8'd21; b = 8'd105;  #10 
a = 8'd21; b = 8'd106;  #10 
a = 8'd21; b = 8'd107;  #10 
a = 8'd21; b = 8'd108;  #10 
a = 8'd21; b = 8'd109;  #10 
a = 8'd21; b = 8'd110;  #10 
a = 8'd21; b = 8'd111;  #10 
a = 8'd21; b = 8'd112;  #10 
a = 8'd21; b = 8'd113;  #10 
a = 8'd21; b = 8'd114;  #10 
a = 8'd21; b = 8'd115;  #10 
a = 8'd21; b = 8'd116;  #10 
a = 8'd21; b = 8'd117;  #10 
a = 8'd21; b = 8'd118;  #10 
a = 8'd21; b = 8'd119;  #10 
a = 8'd21; b = 8'd120;  #10 
a = 8'd21; b = 8'd121;  #10 
a = 8'd21; b = 8'd122;  #10 
a = 8'd21; b = 8'd123;  #10 
a = 8'd21; b = 8'd124;  #10 
a = 8'd21; b = 8'd125;  #10 
a = 8'd21; b = 8'd126;  #10 
a = 8'd21; b = 8'd127;  #10 
a = 8'd21; b = 8'd128;  #10 
a = 8'd21; b = 8'd129;  #10 
a = 8'd21; b = 8'd130;  #10 
a = 8'd21; b = 8'd131;  #10 
a = 8'd21; b = 8'd132;  #10 
a = 8'd21; b = 8'd133;  #10 
a = 8'd21; b = 8'd134;  #10 
a = 8'd21; b = 8'd135;  #10 
a = 8'd21; b = 8'd136;  #10 
a = 8'd21; b = 8'd137;  #10 
a = 8'd21; b = 8'd138;  #10 
a = 8'd21; b = 8'd139;  #10 
a = 8'd21; b = 8'd140;  #10 
a = 8'd21; b = 8'd141;  #10 
a = 8'd21; b = 8'd142;  #10 
a = 8'd21; b = 8'd143;  #10 
a = 8'd21; b = 8'd144;  #10 
a = 8'd21; b = 8'd145;  #10 
a = 8'd21; b = 8'd146;  #10 
a = 8'd21; b = 8'd147;  #10 
a = 8'd21; b = 8'd148;  #10 
a = 8'd21; b = 8'd149;  #10 
a = 8'd21; b = 8'd150;  #10 
a = 8'd21; b = 8'd151;  #10 
a = 8'd21; b = 8'd152;  #10 
a = 8'd21; b = 8'd153;  #10 
a = 8'd21; b = 8'd154;  #10 
a = 8'd21; b = 8'd155;  #10 
a = 8'd21; b = 8'd156;  #10 
a = 8'd21; b = 8'd157;  #10 
a = 8'd21; b = 8'd158;  #10 
a = 8'd21; b = 8'd159;  #10 
a = 8'd21; b = 8'd160;  #10 
a = 8'd21; b = 8'd161;  #10 
a = 8'd21; b = 8'd162;  #10 
a = 8'd21; b = 8'd163;  #10 
a = 8'd21; b = 8'd164;  #10 
a = 8'd21; b = 8'd165;  #10 
a = 8'd21; b = 8'd166;  #10 
a = 8'd21; b = 8'd167;  #10 
a = 8'd21; b = 8'd168;  #10 
a = 8'd21; b = 8'd169;  #10 
a = 8'd21; b = 8'd170;  #10 
a = 8'd21; b = 8'd171;  #10 
a = 8'd21; b = 8'd172;  #10 
a = 8'd21; b = 8'd173;  #10 
a = 8'd21; b = 8'd174;  #10 
a = 8'd21; b = 8'd175;  #10 
a = 8'd21; b = 8'd176;  #10 
a = 8'd21; b = 8'd177;  #10 
a = 8'd21; b = 8'd178;  #10 
a = 8'd21; b = 8'd179;  #10 
a = 8'd21; b = 8'd180;  #10 
a = 8'd21; b = 8'd181;  #10 
a = 8'd21; b = 8'd182;  #10 
a = 8'd21; b = 8'd183;  #10 
a = 8'd21; b = 8'd184;  #10 
a = 8'd21; b = 8'd185;  #10 
a = 8'd21; b = 8'd186;  #10 
a = 8'd21; b = 8'd187;  #10 
a = 8'd21; b = 8'd188;  #10 
a = 8'd21; b = 8'd189;  #10 
a = 8'd21; b = 8'd190;  #10 
a = 8'd21; b = 8'd191;  #10 
a = 8'd21; b = 8'd192;  #10 
a = 8'd21; b = 8'd193;  #10 
a = 8'd21; b = 8'd194;  #10 
a = 8'd21; b = 8'd195;  #10 
a = 8'd21; b = 8'd196;  #10 
a = 8'd21; b = 8'd197;  #10 
a = 8'd21; b = 8'd198;  #10 
a = 8'd21; b = 8'd199;  #10 
a = 8'd21; b = 8'd200;  #10 
a = 8'd21; b = 8'd201;  #10 
a = 8'd21; b = 8'd202;  #10 
a = 8'd21; b = 8'd203;  #10 
a = 8'd21; b = 8'd204;  #10 
a = 8'd21; b = 8'd205;  #10 
a = 8'd21; b = 8'd206;  #10 
a = 8'd21; b = 8'd207;  #10 
a = 8'd21; b = 8'd208;  #10 
a = 8'd21; b = 8'd209;  #10 
a = 8'd21; b = 8'd210;  #10 
a = 8'd21; b = 8'd211;  #10 
a = 8'd21; b = 8'd212;  #10 
a = 8'd21; b = 8'd213;  #10 
a = 8'd21; b = 8'd214;  #10 
a = 8'd21; b = 8'd215;  #10 
a = 8'd21; b = 8'd216;  #10 
a = 8'd21; b = 8'd217;  #10 
a = 8'd21; b = 8'd218;  #10 
a = 8'd21; b = 8'd219;  #10 
a = 8'd21; b = 8'd220;  #10 
a = 8'd21; b = 8'd221;  #10 
a = 8'd21; b = 8'd222;  #10 
a = 8'd21; b = 8'd223;  #10 
a = 8'd21; b = 8'd224;  #10 
a = 8'd21; b = 8'd225;  #10 
a = 8'd21; b = 8'd226;  #10 
a = 8'd21; b = 8'd227;  #10 
a = 8'd21; b = 8'd228;  #10 
a = 8'd21; b = 8'd229;  #10 
a = 8'd21; b = 8'd230;  #10 
a = 8'd21; b = 8'd231;  #10 
a = 8'd21; b = 8'd232;  #10 
a = 8'd21; b = 8'd233;  #10 
a = 8'd21; b = 8'd234;  #10 
a = 8'd21; b = 8'd235;  #10 
a = 8'd21; b = 8'd236;  #10 
a = 8'd21; b = 8'd237;  #10 
a = 8'd21; b = 8'd238;  #10 
a = 8'd21; b = 8'd239;  #10 
a = 8'd21; b = 8'd240;  #10 
a = 8'd21; b = 8'd241;  #10 
a = 8'd21; b = 8'd242;  #10 
a = 8'd21; b = 8'd243;  #10 
a = 8'd21; b = 8'd244;  #10 
a = 8'd21; b = 8'd245;  #10 
a = 8'd21; b = 8'd246;  #10 
a = 8'd21; b = 8'd247;  #10 
a = 8'd21; b = 8'd248;  #10 
a = 8'd21; b = 8'd249;  #10 
a = 8'd21; b = 8'd250;  #10 
a = 8'd21; b = 8'd251;  #10 
a = 8'd21; b = 8'd252;  #10 
a = 8'd21; b = 8'd253;  #10 
a = 8'd21; b = 8'd254;  #10 
a = 8'd21; b = 8'd255;  #10 
a = 8'd22; b = 8'd0;  #10 
a = 8'd22; b = 8'd1;  #10 
a = 8'd22; b = 8'd2;  #10 
a = 8'd22; b = 8'd3;  #10 
a = 8'd22; b = 8'd4;  #10 
a = 8'd22; b = 8'd5;  #10 
a = 8'd22; b = 8'd6;  #10 
a = 8'd22; b = 8'd7;  #10 
a = 8'd22; b = 8'd8;  #10 
a = 8'd22; b = 8'd9;  #10 
a = 8'd22; b = 8'd10;  #10 
a = 8'd22; b = 8'd11;  #10 
a = 8'd22; b = 8'd12;  #10 
a = 8'd22; b = 8'd13;  #10 
a = 8'd22; b = 8'd14;  #10 
a = 8'd22; b = 8'd15;  #10 
a = 8'd22; b = 8'd16;  #10 
a = 8'd22; b = 8'd17;  #10 
a = 8'd22; b = 8'd18;  #10 
a = 8'd22; b = 8'd19;  #10 
a = 8'd22; b = 8'd20;  #10 
a = 8'd22; b = 8'd21;  #10 
a = 8'd22; b = 8'd22;  #10 
a = 8'd22; b = 8'd23;  #10 
a = 8'd22; b = 8'd24;  #10 
a = 8'd22; b = 8'd25;  #10 
a = 8'd22; b = 8'd26;  #10 
a = 8'd22; b = 8'd27;  #10 
a = 8'd22; b = 8'd28;  #10 
a = 8'd22; b = 8'd29;  #10 
a = 8'd22; b = 8'd30;  #10 
a = 8'd22; b = 8'd31;  #10 
a = 8'd22; b = 8'd32;  #10 
a = 8'd22; b = 8'd33;  #10 
a = 8'd22; b = 8'd34;  #10 
a = 8'd22; b = 8'd35;  #10 
a = 8'd22; b = 8'd36;  #10 
a = 8'd22; b = 8'd37;  #10 
a = 8'd22; b = 8'd38;  #10 
a = 8'd22; b = 8'd39;  #10 
a = 8'd22; b = 8'd40;  #10 
a = 8'd22; b = 8'd41;  #10 
a = 8'd22; b = 8'd42;  #10 
a = 8'd22; b = 8'd43;  #10 
a = 8'd22; b = 8'd44;  #10 
a = 8'd22; b = 8'd45;  #10 
a = 8'd22; b = 8'd46;  #10 
a = 8'd22; b = 8'd47;  #10 
a = 8'd22; b = 8'd48;  #10 
a = 8'd22; b = 8'd49;  #10 
a = 8'd22; b = 8'd50;  #10 
a = 8'd22; b = 8'd51;  #10 
a = 8'd22; b = 8'd52;  #10 
a = 8'd22; b = 8'd53;  #10 
a = 8'd22; b = 8'd54;  #10 
a = 8'd22; b = 8'd55;  #10 
a = 8'd22; b = 8'd56;  #10 
a = 8'd22; b = 8'd57;  #10 
a = 8'd22; b = 8'd58;  #10 
a = 8'd22; b = 8'd59;  #10 
a = 8'd22; b = 8'd60;  #10 
a = 8'd22; b = 8'd61;  #10 
a = 8'd22; b = 8'd62;  #10 
a = 8'd22; b = 8'd63;  #10 
a = 8'd22; b = 8'd64;  #10 
a = 8'd22; b = 8'd65;  #10 
a = 8'd22; b = 8'd66;  #10 
a = 8'd22; b = 8'd67;  #10 
a = 8'd22; b = 8'd68;  #10 
a = 8'd22; b = 8'd69;  #10 
a = 8'd22; b = 8'd70;  #10 
a = 8'd22; b = 8'd71;  #10 
a = 8'd22; b = 8'd72;  #10 
a = 8'd22; b = 8'd73;  #10 
a = 8'd22; b = 8'd74;  #10 
a = 8'd22; b = 8'd75;  #10 
a = 8'd22; b = 8'd76;  #10 
a = 8'd22; b = 8'd77;  #10 
a = 8'd22; b = 8'd78;  #10 
a = 8'd22; b = 8'd79;  #10 
a = 8'd22; b = 8'd80;  #10 
a = 8'd22; b = 8'd81;  #10 
a = 8'd22; b = 8'd82;  #10 
a = 8'd22; b = 8'd83;  #10 
a = 8'd22; b = 8'd84;  #10 
a = 8'd22; b = 8'd85;  #10 
a = 8'd22; b = 8'd86;  #10 
a = 8'd22; b = 8'd87;  #10 
a = 8'd22; b = 8'd88;  #10 
a = 8'd22; b = 8'd89;  #10 
a = 8'd22; b = 8'd90;  #10 
a = 8'd22; b = 8'd91;  #10 
a = 8'd22; b = 8'd92;  #10 
a = 8'd22; b = 8'd93;  #10 
a = 8'd22; b = 8'd94;  #10 
a = 8'd22; b = 8'd95;  #10 
a = 8'd22; b = 8'd96;  #10 
a = 8'd22; b = 8'd97;  #10 
a = 8'd22; b = 8'd98;  #10 
a = 8'd22; b = 8'd99;  #10 
a = 8'd22; b = 8'd100;  #10 
a = 8'd22; b = 8'd101;  #10 
a = 8'd22; b = 8'd102;  #10 
a = 8'd22; b = 8'd103;  #10 
a = 8'd22; b = 8'd104;  #10 
a = 8'd22; b = 8'd105;  #10 
a = 8'd22; b = 8'd106;  #10 
a = 8'd22; b = 8'd107;  #10 
a = 8'd22; b = 8'd108;  #10 
a = 8'd22; b = 8'd109;  #10 
a = 8'd22; b = 8'd110;  #10 
a = 8'd22; b = 8'd111;  #10 
a = 8'd22; b = 8'd112;  #10 
a = 8'd22; b = 8'd113;  #10 
a = 8'd22; b = 8'd114;  #10 
a = 8'd22; b = 8'd115;  #10 
a = 8'd22; b = 8'd116;  #10 
a = 8'd22; b = 8'd117;  #10 
a = 8'd22; b = 8'd118;  #10 
a = 8'd22; b = 8'd119;  #10 
a = 8'd22; b = 8'd120;  #10 
a = 8'd22; b = 8'd121;  #10 
a = 8'd22; b = 8'd122;  #10 
a = 8'd22; b = 8'd123;  #10 
a = 8'd22; b = 8'd124;  #10 
a = 8'd22; b = 8'd125;  #10 
a = 8'd22; b = 8'd126;  #10 
a = 8'd22; b = 8'd127;  #10 
a = 8'd22; b = 8'd128;  #10 
a = 8'd22; b = 8'd129;  #10 
a = 8'd22; b = 8'd130;  #10 
a = 8'd22; b = 8'd131;  #10 
a = 8'd22; b = 8'd132;  #10 
a = 8'd22; b = 8'd133;  #10 
a = 8'd22; b = 8'd134;  #10 
a = 8'd22; b = 8'd135;  #10 
a = 8'd22; b = 8'd136;  #10 
a = 8'd22; b = 8'd137;  #10 
a = 8'd22; b = 8'd138;  #10 
a = 8'd22; b = 8'd139;  #10 
a = 8'd22; b = 8'd140;  #10 
a = 8'd22; b = 8'd141;  #10 
a = 8'd22; b = 8'd142;  #10 
a = 8'd22; b = 8'd143;  #10 
a = 8'd22; b = 8'd144;  #10 
a = 8'd22; b = 8'd145;  #10 
a = 8'd22; b = 8'd146;  #10 
a = 8'd22; b = 8'd147;  #10 
a = 8'd22; b = 8'd148;  #10 
a = 8'd22; b = 8'd149;  #10 
a = 8'd22; b = 8'd150;  #10 
a = 8'd22; b = 8'd151;  #10 
a = 8'd22; b = 8'd152;  #10 
a = 8'd22; b = 8'd153;  #10 
a = 8'd22; b = 8'd154;  #10 
a = 8'd22; b = 8'd155;  #10 
a = 8'd22; b = 8'd156;  #10 
a = 8'd22; b = 8'd157;  #10 
a = 8'd22; b = 8'd158;  #10 
a = 8'd22; b = 8'd159;  #10 
a = 8'd22; b = 8'd160;  #10 
a = 8'd22; b = 8'd161;  #10 
a = 8'd22; b = 8'd162;  #10 
a = 8'd22; b = 8'd163;  #10 
a = 8'd22; b = 8'd164;  #10 
a = 8'd22; b = 8'd165;  #10 
a = 8'd22; b = 8'd166;  #10 
a = 8'd22; b = 8'd167;  #10 
a = 8'd22; b = 8'd168;  #10 
a = 8'd22; b = 8'd169;  #10 
a = 8'd22; b = 8'd170;  #10 
a = 8'd22; b = 8'd171;  #10 
a = 8'd22; b = 8'd172;  #10 
a = 8'd22; b = 8'd173;  #10 
a = 8'd22; b = 8'd174;  #10 
a = 8'd22; b = 8'd175;  #10 
a = 8'd22; b = 8'd176;  #10 
a = 8'd22; b = 8'd177;  #10 
a = 8'd22; b = 8'd178;  #10 
a = 8'd22; b = 8'd179;  #10 
a = 8'd22; b = 8'd180;  #10 
a = 8'd22; b = 8'd181;  #10 
a = 8'd22; b = 8'd182;  #10 
a = 8'd22; b = 8'd183;  #10 
a = 8'd22; b = 8'd184;  #10 
a = 8'd22; b = 8'd185;  #10 
a = 8'd22; b = 8'd186;  #10 
a = 8'd22; b = 8'd187;  #10 
a = 8'd22; b = 8'd188;  #10 
a = 8'd22; b = 8'd189;  #10 
a = 8'd22; b = 8'd190;  #10 
a = 8'd22; b = 8'd191;  #10 
a = 8'd22; b = 8'd192;  #10 
a = 8'd22; b = 8'd193;  #10 
a = 8'd22; b = 8'd194;  #10 
a = 8'd22; b = 8'd195;  #10 
a = 8'd22; b = 8'd196;  #10 
a = 8'd22; b = 8'd197;  #10 
a = 8'd22; b = 8'd198;  #10 
a = 8'd22; b = 8'd199;  #10 
a = 8'd22; b = 8'd200;  #10 
a = 8'd22; b = 8'd201;  #10 
a = 8'd22; b = 8'd202;  #10 
a = 8'd22; b = 8'd203;  #10 
a = 8'd22; b = 8'd204;  #10 
a = 8'd22; b = 8'd205;  #10 
a = 8'd22; b = 8'd206;  #10 
a = 8'd22; b = 8'd207;  #10 
a = 8'd22; b = 8'd208;  #10 
a = 8'd22; b = 8'd209;  #10 
a = 8'd22; b = 8'd210;  #10 
a = 8'd22; b = 8'd211;  #10 
a = 8'd22; b = 8'd212;  #10 
a = 8'd22; b = 8'd213;  #10 
a = 8'd22; b = 8'd214;  #10 
a = 8'd22; b = 8'd215;  #10 
a = 8'd22; b = 8'd216;  #10 
a = 8'd22; b = 8'd217;  #10 
a = 8'd22; b = 8'd218;  #10 
a = 8'd22; b = 8'd219;  #10 
a = 8'd22; b = 8'd220;  #10 
a = 8'd22; b = 8'd221;  #10 
a = 8'd22; b = 8'd222;  #10 
a = 8'd22; b = 8'd223;  #10 
a = 8'd22; b = 8'd224;  #10 
a = 8'd22; b = 8'd225;  #10 
a = 8'd22; b = 8'd226;  #10 
a = 8'd22; b = 8'd227;  #10 
a = 8'd22; b = 8'd228;  #10 
a = 8'd22; b = 8'd229;  #10 
a = 8'd22; b = 8'd230;  #10 
a = 8'd22; b = 8'd231;  #10 
a = 8'd22; b = 8'd232;  #10 
a = 8'd22; b = 8'd233;  #10 
a = 8'd22; b = 8'd234;  #10 
a = 8'd22; b = 8'd235;  #10 
a = 8'd22; b = 8'd236;  #10 
a = 8'd22; b = 8'd237;  #10 
a = 8'd22; b = 8'd238;  #10 
a = 8'd22; b = 8'd239;  #10 
a = 8'd22; b = 8'd240;  #10 
a = 8'd22; b = 8'd241;  #10 
a = 8'd22; b = 8'd242;  #10 
a = 8'd22; b = 8'd243;  #10 
a = 8'd22; b = 8'd244;  #10 
a = 8'd22; b = 8'd245;  #10 
a = 8'd22; b = 8'd246;  #10 
a = 8'd22; b = 8'd247;  #10 
a = 8'd22; b = 8'd248;  #10 
a = 8'd22; b = 8'd249;  #10 
a = 8'd22; b = 8'd250;  #10 
a = 8'd22; b = 8'd251;  #10 
a = 8'd22; b = 8'd252;  #10 
a = 8'd22; b = 8'd253;  #10 
a = 8'd22; b = 8'd254;  #10 
a = 8'd22; b = 8'd255;  #10 
a = 8'd23; b = 8'd0;  #10 
a = 8'd23; b = 8'd1;  #10 
a = 8'd23; b = 8'd2;  #10 
a = 8'd23; b = 8'd3;  #10 
a = 8'd23; b = 8'd4;  #10 
a = 8'd23; b = 8'd5;  #10 
a = 8'd23; b = 8'd6;  #10 
a = 8'd23; b = 8'd7;  #10 
a = 8'd23; b = 8'd8;  #10 
a = 8'd23; b = 8'd9;  #10 
a = 8'd23; b = 8'd10;  #10 
a = 8'd23; b = 8'd11;  #10 
a = 8'd23; b = 8'd12;  #10 
a = 8'd23; b = 8'd13;  #10 
a = 8'd23; b = 8'd14;  #10 
a = 8'd23; b = 8'd15;  #10 
a = 8'd23; b = 8'd16;  #10 
a = 8'd23; b = 8'd17;  #10 
a = 8'd23; b = 8'd18;  #10 
a = 8'd23; b = 8'd19;  #10 
a = 8'd23; b = 8'd20;  #10 
a = 8'd23; b = 8'd21;  #10 
a = 8'd23; b = 8'd22;  #10 
a = 8'd23; b = 8'd23;  #10 
a = 8'd23; b = 8'd24;  #10 
a = 8'd23; b = 8'd25;  #10 
a = 8'd23; b = 8'd26;  #10 
a = 8'd23; b = 8'd27;  #10 
a = 8'd23; b = 8'd28;  #10 
a = 8'd23; b = 8'd29;  #10 
a = 8'd23; b = 8'd30;  #10 
a = 8'd23; b = 8'd31;  #10 
a = 8'd23; b = 8'd32;  #10 
a = 8'd23; b = 8'd33;  #10 
a = 8'd23; b = 8'd34;  #10 
a = 8'd23; b = 8'd35;  #10 
a = 8'd23; b = 8'd36;  #10 
a = 8'd23; b = 8'd37;  #10 
a = 8'd23; b = 8'd38;  #10 
a = 8'd23; b = 8'd39;  #10 
a = 8'd23; b = 8'd40;  #10 
a = 8'd23; b = 8'd41;  #10 
a = 8'd23; b = 8'd42;  #10 
a = 8'd23; b = 8'd43;  #10 
a = 8'd23; b = 8'd44;  #10 
a = 8'd23; b = 8'd45;  #10 
a = 8'd23; b = 8'd46;  #10 
a = 8'd23; b = 8'd47;  #10 
a = 8'd23; b = 8'd48;  #10 
a = 8'd23; b = 8'd49;  #10 
a = 8'd23; b = 8'd50;  #10 
a = 8'd23; b = 8'd51;  #10 
a = 8'd23; b = 8'd52;  #10 
a = 8'd23; b = 8'd53;  #10 
a = 8'd23; b = 8'd54;  #10 
a = 8'd23; b = 8'd55;  #10 
a = 8'd23; b = 8'd56;  #10 
a = 8'd23; b = 8'd57;  #10 
a = 8'd23; b = 8'd58;  #10 
a = 8'd23; b = 8'd59;  #10 
a = 8'd23; b = 8'd60;  #10 
a = 8'd23; b = 8'd61;  #10 
a = 8'd23; b = 8'd62;  #10 
a = 8'd23; b = 8'd63;  #10 
a = 8'd23; b = 8'd64;  #10 
a = 8'd23; b = 8'd65;  #10 
a = 8'd23; b = 8'd66;  #10 
a = 8'd23; b = 8'd67;  #10 
a = 8'd23; b = 8'd68;  #10 
a = 8'd23; b = 8'd69;  #10 
a = 8'd23; b = 8'd70;  #10 
a = 8'd23; b = 8'd71;  #10 
a = 8'd23; b = 8'd72;  #10 
a = 8'd23; b = 8'd73;  #10 
a = 8'd23; b = 8'd74;  #10 
a = 8'd23; b = 8'd75;  #10 
a = 8'd23; b = 8'd76;  #10 
a = 8'd23; b = 8'd77;  #10 
a = 8'd23; b = 8'd78;  #10 
a = 8'd23; b = 8'd79;  #10 
a = 8'd23; b = 8'd80;  #10 
a = 8'd23; b = 8'd81;  #10 
a = 8'd23; b = 8'd82;  #10 
a = 8'd23; b = 8'd83;  #10 
a = 8'd23; b = 8'd84;  #10 
a = 8'd23; b = 8'd85;  #10 
a = 8'd23; b = 8'd86;  #10 
a = 8'd23; b = 8'd87;  #10 
a = 8'd23; b = 8'd88;  #10 
a = 8'd23; b = 8'd89;  #10 
a = 8'd23; b = 8'd90;  #10 
a = 8'd23; b = 8'd91;  #10 
a = 8'd23; b = 8'd92;  #10 
a = 8'd23; b = 8'd93;  #10 
a = 8'd23; b = 8'd94;  #10 
a = 8'd23; b = 8'd95;  #10 
a = 8'd23; b = 8'd96;  #10 
a = 8'd23; b = 8'd97;  #10 
a = 8'd23; b = 8'd98;  #10 
a = 8'd23; b = 8'd99;  #10 
a = 8'd23; b = 8'd100;  #10 
a = 8'd23; b = 8'd101;  #10 
a = 8'd23; b = 8'd102;  #10 
a = 8'd23; b = 8'd103;  #10 
a = 8'd23; b = 8'd104;  #10 
a = 8'd23; b = 8'd105;  #10 
a = 8'd23; b = 8'd106;  #10 
a = 8'd23; b = 8'd107;  #10 
a = 8'd23; b = 8'd108;  #10 
a = 8'd23; b = 8'd109;  #10 
a = 8'd23; b = 8'd110;  #10 
a = 8'd23; b = 8'd111;  #10 
a = 8'd23; b = 8'd112;  #10 
a = 8'd23; b = 8'd113;  #10 
a = 8'd23; b = 8'd114;  #10 
a = 8'd23; b = 8'd115;  #10 
a = 8'd23; b = 8'd116;  #10 
a = 8'd23; b = 8'd117;  #10 
a = 8'd23; b = 8'd118;  #10 
a = 8'd23; b = 8'd119;  #10 
a = 8'd23; b = 8'd120;  #10 
a = 8'd23; b = 8'd121;  #10 
a = 8'd23; b = 8'd122;  #10 
a = 8'd23; b = 8'd123;  #10 
a = 8'd23; b = 8'd124;  #10 
a = 8'd23; b = 8'd125;  #10 
a = 8'd23; b = 8'd126;  #10 
a = 8'd23; b = 8'd127;  #10 
a = 8'd23; b = 8'd128;  #10 
a = 8'd23; b = 8'd129;  #10 
a = 8'd23; b = 8'd130;  #10 
a = 8'd23; b = 8'd131;  #10 
a = 8'd23; b = 8'd132;  #10 
a = 8'd23; b = 8'd133;  #10 
a = 8'd23; b = 8'd134;  #10 
a = 8'd23; b = 8'd135;  #10 
a = 8'd23; b = 8'd136;  #10 
a = 8'd23; b = 8'd137;  #10 
a = 8'd23; b = 8'd138;  #10 
a = 8'd23; b = 8'd139;  #10 
a = 8'd23; b = 8'd140;  #10 
a = 8'd23; b = 8'd141;  #10 
a = 8'd23; b = 8'd142;  #10 
a = 8'd23; b = 8'd143;  #10 
a = 8'd23; b = 8'd144;  #10 
a = 8'd23; b = 8'd145;  #10 
a = 8'd23; b = 8'd146;  #10 
a = 8'd23; b = 8'd147;  #10 
a = 8'd23; b = 8'd148;  #10 
a = 8'd23; b = 8'd149;  #10 
a = 8'd23; b = 8'd150;  #10 
a = 8'd23; b = 8'd151;  #10 
a = 8'd23; b = 8'd152;  #10 
a = 8'd23; b = 8'd153;  #10 
a = 8'd23; b = 8'd154;  #10 
a = 8'd23; b = 8'd155;  #10 
a = 8'd23; b = 8'd156;  #10 
a = 8'd23; b = 8'd157;  #10 
a = 8'd23; b = 8'd158;  #10 
a = 8'd23; b = 8'd159;  #10 
a = 8'd23; b = 8'd160;  #10 
a = 8'd23; b = 8'd161;  #10 
a = 8'd23; b = 8'd162;  #10 
a = 8'd23; b = 8'd163;  #10 
a = 8'd23; b = 8'd164;  #10 
a = 8'd23; b = 8'd165;  #10 
a = 8'd23; b = 8'd166;  #10 
a = 8'd23; b = 8'd167;  #10 
a = 8'd23; b = 8'd168;  #10 
a = 8'd23; b = 8'd169;  #10 
a = 8'd23; b = 8'd170;  #10 
a = 8'd23; b = 8'd171;  #10 
a = 8'd23; b = 8'd172;  #10 
a = 8'd23; b = 8'd173;  #10 
a = 8'd23; b = 8'd174;  #10 
a = 8'd23; b = 8'd175;  #10 
a = 8'd23; b = 8'd176;  #10 
a = 8'd23; b = 8'd177;  #10 
a = 8'd23; b = 8'd178;  #10 
a = 8'd23; b = 8'd179;  #10 
a = 8'd23; b = 8'd180;  #10 
a = 8'd23; b = 8'd181;  #10 
a = 8'd23; b = 8'd182;  #10 
a = 8'd23; b = 8'd183;  #10 
a = 8'd23; b = 8'd184;  #10 
a = 8'd23; b = 8'd185;  #10 
a = 8'd23; b = 8'd186;  #10 
a = 8'd23; b = 8'd187;  #10 
a = 8'd23; b = 8'd188;  #10 
a = 8'd23; b = 8'd189;  #10 
a = 8'd23; b = 8'd190;  #10 
a = 8'd23; b = 8'd191;  #10 
a = 8'd23; b = 8'd192;  #10 
a = 8'd23; b = 8'd193;  #10 
a = 8'd23; b = 8'd194;  #10 
a = 8'd23; b = 8'd195;  #10 
a = 8'd23; b = 8'd196;  #10 
a = 8'd23; b = 8'd197;  #10 
a = 8'd23; b = 8'd198;  #10 
a = 8'd23; b = 8'd199;  #10 
a = 8'd23; b = 8'd200;  #10 
a = 8'd23; b = 8'd201;  #10 
a = 8'd23; b = 8'd202;  #10 
a = 8'd23; b = 8'd203;  #10 
a = 8'd23; b = 8'd204;  #10 
a = 8'd23; b = 8'd205;  #10 
a = 8'd23; b = 8'd206;  #10 
a = 8'd23; b = 8'd207;  #10 
a = 8'd23; b = 8'd208;  #10 
a = 8'd23; b = 8'd209;  #10 
a = 8'd23; b = 8'd210;  #10 
a = 8'd23; b = 8'd211;  #10 
a = 8'd23; b = 8'd212;  #10 
a = 8'd23; b = 8'd213;  #10 
a = 8'd23; b = 8'd214;  #10 
a = 8'd23; b = 8'd215;  #10 
a = 8'd23; b = 8'd216;  #10 
a = 8'd23; b = 8'd217;  #10 
a = 8'd23; b = 8'd218;  #10 
a = 8'd23; b = 8'd219;  #10 
a = 8'd23; b = 8'd220;  #10 
a = 8'd23; b = 8'd221;  #10 
a = 8'd23; b = 8'd222;  #10 
a = 8'd23; b = 8'd223;  #10 
a = 8'd23; b = 8'd224;  #10 
a = 8'd23; b = 8'd225;  #10 
a = 8'd23; b = 8'd226;  #10 
a = 8'd23; b = 8'd227;  #10 
a = 8'd23; b = 8'd228;  #10 
a = 8'd23; b = 8'd229;  #10 
a = 8'd23; b = 8'd230;  #10 
a = 8'd23; b = 8'd231;  #10 
a = 8'd23; b = 8'd232;  #10 
a = 8'd23; b = 8'd233;  #10 
a = 8'd23; b = 8'd234;  #10 
a = 8'd23; b = 8'd235;  #10 
a = 8'd23; b = 8'd236;  #10 
a = 8'd23; b = 8'd237;  #10 
a = 8'd23; b = 8'd238;  #10 
a = 8'd23; b = 8'd239;  #10 
a = 8'd23; b = 8'd240;  #10 
a = 8'd23; b = 8'd241;  #10 
a = 8'd23; b = 8'd242;  #10 
a = 8'd23; b = 8'd243;  #10 
a = 8'd23; b = 8'd244;  #10 
a = 8'd23; b = 8'd245;  #10 
a = 8'd23; b = 8'd246;  #10 
a = 8'd23; b = 8'd247;  #10 
a = 8'd23; b = 8'd248;  #10 
a = 8'd23; b = 8'd249;  #10 
a = 8'd23; b = 8'd250;  #10 
a = 8'd23; b = 8'd251;  #10 
a = 8'd23; b = 8'd252;  #10 
a = 8'd23; b = 8'd253;  #10 
a = 8'd23; b = 8'd254;  #10 
a = 8'd23; b = 8'd255;  #10 
a = 8'd24; b = 8'd0;  #10 
a = 8'd24; b = 8'd1;  #10 
a = 8'd24; b = 8'd2;  #10 
a = 8'd24; b = 8'd3;  #10 
a = 8'd24; b = 8'd4;  #10 
a = 8'd24; b = 8'd5;  #10 
a = 8'd24; b = 8'd6;  #10 
a = 8'd24; b = 8'd7;  #10 
a = 8'd24; b = 8'd8;  #10 
a = 8'd24; b = 8'd9;  #10 
a = 8'd24; b = 8'd10;  #10 
a = 8'd24; b = 8'd11;  #10 
a = 8'd24; b = 8'd12;  #10 
a = 8'd24; b = 8'd13;  #10 
a = 8'd24; b = 8'd14;  #10 
a = 8'd24; b = 8'd15;  #10 
a = 8'd24; b = 8'd16;  #10 
a = 8'd24; b = 8'd17;  #10 
a = 8'd24; b = 8'd18;  #10 
a = 8'd24; b = 8'd19;  #10 
a = 8'd24; b = 8'd20;  #10 
a = 8'd24; b = 8'd21;  #10 
a = 8'd24; b = 8'd22;  #10 
a = 8'd24; b = 8'd23;  #10 
a = 8'd24; b = 8'd24;  #10 
a = 8'd24; b = 8'd25;  #10 
a = 8'd24; b = 8'd26;  #10 
a = 8'd24; b = 8'd27;  #10 
a = 8'd24; b = 8'd28;  #10 
a = 8'd24; b = 8'd29;  #10 
a = 8'd24; b = 8'd30;  #10 
a = 8'd24; b = 8'd31;  #10 
a = 8'd24; b = 8'd32;  #10 
a = 8'd24; b = 8'd33;  #10 
a = 8'd24; b = 8'd34;  #10 
a = 8'd24; b = 8'd35;  #10 
a = 8'd24; b = 8'd36;  #10 
a = 8'd24; b = 8'd37;  #10 
a = 8'd24; b = 8'd38;  #10 
a = 8'd24; b = 8'd39;  #10 
a = 8'd24; b = 8'd40;  #10 
a = 8'd24; b = 8'd41;  #10 
a = 8'd24; b = 8'd42;  #10 
a = 8'd24; b = 8'd43;  #10 
a = 8'd24; b = 8'd44;  #10 
a = 8'd24; b = 8'd45;  #10 
a = 8'd24; b = 8'd46;  #10 
a = 8'd24; b = 8'd47;  #10 
a = 8'd24; b = 8'd48;  #10 
a = 8'd24; b = 8'd49;  #10 
a = 8'd24; b = 8'd50;  #10 
a = 8'd24; b = 8'd51;  #10 
a = 8'd24; b = 8'd52;  #10 
a = 8'd24; b = 8'd53;  #10 
a = 8'd24; b = 8'd54;  #10 
a = 8'd24; b = 8'd55;  #10 
a = 8'd24; b = 8'd56;  #10 
a = 8'd24; b = 8'd57;  #10 
a = 8'd24; b = 8'd58;  #10 
a = 8'd24; b = 8'd59;  #10 
a = 8'd24; b = 8'd60;  #10 
a = 8'd24; b = 8'd61;  #10 
a = 8'd24; b = 8'd62;  #10 
a = 8'd24; b = 8'd63;  #10 
a = 8'd24; b = 8'd64;  #10 
a = 8'd24; b = 8'd65;  #10 
a = 8'd24; b = 8'd66;  #10 
a = 8'd24; b = 8'd67;  #10 
a = 8'd24; b = 8'd68;  #10 
a = 8'd24; b = 8'd69;  #10 
a = 8'd24; b = 8'd70;  #10 
a = 8'd24; b = 8'd71;  #10 
a = 8'd24; b = 8'd72;  #10 
a = 8'd24; b = 8'd73;  #10 
a = 8'd24; b = 8'd74;  #10 
a = 8'd24; b = 8'd75;  #10 
a = 8'd24; b = 8'd76;  #10 
a = 8'd24; b = 8'd77;  #10 
a = 8'd24; b = 8'd78;  #10 
a = 8'd24; b = 8'd79;  #10 
a = 8'd24; b = 8'd80;  #10 
a = 8'd24; b = 8'd81;  #10 
a = 8'd24; b = 8'd82;  #10 
a = 8'd24; b = 8'd83;  #10 
a = 8'd24; b = 8'd84;  #10 
a = 8'd24; b = 8'd85;  #10 
a = 8'd24; b = 8'd86;  #10 
a = 8'd24; b = 8'd87;  #10 
a = 8'd24; b = 8'd88;  #10 
a = 8'd24; b = 8'd89;  #10 
a = 8'd24; b = 8'd90;  #10 
a = 8'd24; b = 8'd91;  #10 
a = 8'd24; b = 8'd92;  #10 
a = 8'd24; b = 8'd93;  #10 
a = 8'd24; b = 8'd94;  #10 
a = 8'd24; b = 8'd95;  #10 
a = 8'd24; b = 8'd96;  #10 
a = 8'd24; b = 8'd97;  #10 
a = 8'd24; b = 8'd98;  #10 
a = 8'd24; b = 8'd99;  #10 
a = 8'd24; b = 8'd100;  #10 
a = 8'd24; b = 8'd101;  #10 
a = 8'd24; b = 8'd102;  #10 
a = 8'd24; b = 8'd103;  #10 
a = 8'd24; b = 8'd104;  #10 
a = 8'd24; b = 8'd105;  #10 
a = 8'd24; b = 8'd106;  #10 
a = 8'd24; b = 8'd107;  #10 
a = 8'd24; b = 8'd108;  #10 
a = 8'd24; b = 8'd109;  #10 
a = 8'd24; b = 8'd110;  #10 
a = 8'd24; b = 8'd111;  #10 
a = 8'd24; b = 8'd112;  #10 
a = 8'd24; b = 8'd113;  #10 
a = 8'd24; b = 8'd114;  #10 
a = 8'd24; b = 8'd115;  #10 
a = 8'd24; b = 8'd116;  #10 
a = 8'd24; b = 8'd117;  #10 
a = 8'd24; b = 8'd118;  #10 
a = 8'd24; b = 8'd119;  #10 
a = 8'd24; b = 8'd120;  #10 
a = 8'd24; b = 8'd121;  #10 
a = 8'd24; b = 8'd122;  #10 
a = 8'd24; b = 8'd123;  #10 
a = 8'd24; b = 8'd124;  #10 
a = 8'd24; b = 8'd125;  #10 
a = 8'd24; b = 8'd126;  #10 
a = 8'd24; b = 8'd127;  #10 
a = 8'd24; b = 8'd128;  #10 
a = 8'd24; b = 8'd129;  #10 
a = 8'd24; b = 8'd130;  #10 
a = 8'd24; b = 8'd131;  #10 
a = 8'd24; b = 8'd132;  #10 
a = 8'd24; b = 8'd133;  #10 
a = 8'd24; b = 8'd134;  #10 
a = 8'd24; b = 8'd135;  #10 
a = 8'd24; b = 8'd136;  #10 
a = 8'd24; b = 8'd137;  #10 
a = 8'd24; b = 8'd138;  #10 
a = 8'd24; b = 8'd139;  #10 
a = 8'd24; b = 8'd140;  #10 
a = 8'd24; b = 8'd141;  #10 
a = 8'd24; b = 8'd142;  #10 
a = 8'd24; b = 8'd143;  #10 
a = 8'd24; b = 8'd144;  #10 
a = 8'd24; b = 8'd145;  #10 
a = 8'd24; b = 8'd146;  #10 
a = 8'd24; b = 8'd147;  #10 
a = 8'd24; b = 8'd148;  #10 
a = 8'd24; b = 8'd149;  #10 
a = 8'd24; b = 8'd150;  #10 
a = 8'd24; b = 8'd151;  #10 
a = 8'd24; b = 8'd152;  #10 
a = 8'd24; b = 8'd153;  #10 
a = 8'd24; b = 8'd154;  #10 
a = 8'd24; b = 8'd155;  #10 
a = 8'd24; b = 8'd156;  #10 
a = 8'd24; b = 8'd157;  #10 
a = 8'd24; b = 8'd158;  #10 
a = 8'd24; b = 8'd159;  #10 
a = 8'd24; b = 8'd160;  #10 
a = 8'd24; b = 8'd161;  #10 
a = 8'd24; b = 8'd162;  #10 
a = 8'd24; b = 8'd163;  #10 
a = 8'd24; b = 8'd164;  #10 
a = 8'd24; b = 8'd165;  #10 
a = 8'd24; b = 8'd166;  #10 
a = 8'd24; b = 8'd167;  #10 
a = 8'd24; b = 8'd168;  #10 
a = 8'd24; b = 8'd169;  #10 
a = 8'd24; b = 8'd170;  #10 
a = 8'd24; b = 8'd171;  #10 
a = 8'd24; b = 8'd172;  #10 
a = 8'd24; b = 8'd173;  #10 
a = 8'd24; b = 8'd174;  #10 
a = 8'd24; b = 8'd175;  #10 
a = 8'd24; b = 8'd176;  #10 
a = 8'd24; b = 8'd177;  #10 
a = 8'd24; b = 8'd178;  #10 
a = 8'd24; b = 8'd179;  #10 
a = 8'd24; b = 8'd180;  #10 
a = 8'd24; b = 8'd181;  #10 
a = 8'd24; b = 8'd182;  #10 
a = 8'd24; b = 8'd183;  #10 
a = 8'd24; b = 8'd184;  #10 
a = 8'd24; b = 8'd185;  #10 
a = 8'd24; b = 8'd186;  #10 
a = 8'd24; b = 8'd187;  #10 
a = 8'd24; b = 8'd188;  #10 
a = 8'd24; b = 8'd189;  #10 
a = 8'd24; b = 8'd190;  #10 
a = 8'd24; b = 8'd191;  #10 
a = 8'd24; b = 8'd192;  #10 
a = 8'd24; b = 8'd193;  #10 
a = 8'd24; b = 8'd194;  #10 
a = 8'd24; b = 8'd195;  #10 
a = 8'd24; b = 8'd196;  #10 
a = 8'd24; b = 8'd197;  #10 
a = 8'd24; b = 8'd198;  #10 
a = 8'd24; b = 8'd199;  #10 
a = 8'd24; b = 8'd200;  #10 
a = 8'd24; b = 8'd201;  #10 
a = 8'd24; b = 8'd202;  #10 
a = 8'd24; b = 8'd203;  #10 
a = 8'd24; b = 8'd204;  #10 
a = 8'd24; b = 8'd205;  #10 
a = 8'd24; b = 8'd206;  #10 
a = 8'd24; b = 8'd207;  #10 
a = 8'd24; b = 8'd208;  #10 
a = 8'd24; b = 8'd209;  #10 
a = 8'd24; b = 8'd210;  #10 
a = 8'd24; b = 8'd211;  #10 
a = 8'd24; b = 8'd212;  #10 
a = 8'd24; b = 8'd213;  #10 
a = 8'd24; b = 8'd214;  #10 
a = 8'd24; b = 8'd215;  #10 
a = 8'd24; b = 8'd216;  #10 
a = 8'd24; b = 8'd217;  #10 
a = 8'd24; b = 8'd218;  #10 
a = 8'd24; b = 8'd219;  #10 
a = 8'd24; b = 8'd220;  #10 
a = 8'd24; b = 8'd221;  #10 
a = 8'd24; b = 8'd222;  #10 
a = 8'd24; b = 8'd223;  #10 
a = 8'd24; b = 8'd224;  #10 
a = 8'd24; b = 8'd225;  #10 
a = 8'd24; b = 8'd226;  #10 
a = 8'd24; b = 8'd227;  #10 
a = 8'd24; b = 8'd228;  #10 
a = 8'd24; b = 8'd229;  #10 
a = 8'd24; b = 8'd230;  #10 
a = 8'd24; b = 8'd231;  #10 
a = 8'd24; b = 8'd232;  #10 
a = 8'd24; b = 8'd233;  #10 
a = 8'd24; b = 8'd234;  #10 
a = 8'd24; b = 8'd235;  #10 
a = 8'd24; b = 8'd236;  #10 
a = 8'd24; b = 8'd237;  #10 
a = 8'd24; b = 8'd238;  #10 
a = 8'd24; b = 8'd239;  #10 
a = 8'd24; b = 8'd240;  #10 
a = 8'd24; b = 8'd241;  #10 
a = 8'd24; b = 8'd242;  #10 
a = 8'd24; b = 8'd243;  #10 
a = 8'd24; b = 8'd244;  #10 
a = 8'd24; b = 8'd245;  #10 
a = 8'd24; b = 8'd246;  #10 
a = 8'd24; b = 8'd247;  #10 
a = 8'd24; b = 8'd248;  #10 
a = 8'd24; b = 8'd249;  #10 
a = 8'd24; b = 8'd250;  #10 
a = 8'd24; b = 8'd251;  #10 
a = 8'd24; b = 8'd252;  #10 
a = 8'd24; b = 8'd253;  #10 
a = 8'd24; b = 8'd254;  #10 
a = 8'd24; b = 8'd255;  #10 
a = 8'd25; b = 8'd0;  #10 
a = 8'd25; b = 8'd1;  #10 
a = 8'd25; b = 8'd2;  #10 
a = 8'd25; b = 8'd3;  #10 
a = 8'd25; b = 8'd4;  #10 
a = 8'd25; b = 8'd5;  #10 
a = 8'd25; b = 8'd6;  #10 
a = 8'd25; b = 8'd7;  #10 
a = 8'd25; b = 8'd8;  #10 
a = 8'd25; b = 8'd9;  #10 
a = 8'd25; b = 8'd10;  #10 
a = 8'd25; b = 8'd11;  #10 
a = 8'd25; b = 8'd12;  #10 
a = 8'd25; b = 8'd13;  #10 
a = 8'd25; b = 8'd14;  #10 
a = 8'd25; b = 8'd15;  #10 
a = 8'd25; b = 8'd16;  #10 
a = 8'd25; b = 8'd17;  #10 
a = 8'd25; b = 8'd18;  #10 
a = 8'd25; b = 8'd19;  #10 
a = 8'd25; b = 8'd20;  #10 
a = 8'd25; b = 8'd21;  #10 
a = 8'd25; b = 8'd22;  #10 
a = 8'd25; b = 8'd23;  #10 
a = 8'd25; b = 8'd24;  #10 
a = 8'd25; b = 8'd25;  #10 
a = 8'd25; b = 8'd26;  #10 
a = 8'd25; b = 8'd27;  #10 
a = 8'd25; b = 8'd28;  #10 
a = 8'd25; b = 8'd29;  #10 
a = 8'd25; b = 8'd30;  #10 
a = 8'd25; b = 8'd31;  #10 
a = 8'd25; b = 8'd32;  #10 
a = 8'd25; b = 8'd33;  #10 
a = 8'd25; b = 8'd34;  #10 
a = 8'd25; b = 8'd35;  #10 
a = 8'd25; b = 8'd36;  #10 
a = 8'd25; b = 8'd37;  #10 
a = 8'd25; b = 8'd38;  #10 
a = 8'd25; b = 8'd39;  #10 
a = 8'd25; b = 8'd40;  #10 
a = 8'd25; b = 8'd41;  #10 
a = 8'd25; b = 8'd42;  #10 
a = 8'd25; b = 8'd43;  #10 
a = 8'd25; b = 8'd44;  #10 
a = 8'd25; b = 8'd45;  #10 
a = 8'd25; b = 8'd46;  #10 
a = 8'd25; b = 8'd47;  #10 
a = 8'd25; b = 8'd48;  #10 
a = 8'd25; b = 8'd49;  #10 
a = 8'd25; b = 8'd50;  #10 
a = 8'd25; b = 8'd51;  #10 
a = 8'd25; b = 8'd52;  #10 
a = 8'd25; b = 8'd53;  #10 
a = 8'd25; b = 8'd54;  #10 
a = 8'd25; b = 8'd55;  #10 
a = 8'd25; b = 8'd56;  #10 
a = 8'd25; b = 8'd57;  #10 
a = 8'd25; b = 8'd58;  #10 
a = 8'd25; b = 8'd59;  #10 
a = 8'd25; b = 8'd60;  #10 
a = 8'd25; b = 8'd61;  #10 
a = 8'd25; b = 8'd62;  #10 
a = 8'd25; b = 8'd63;  #10 
a = 8'd25; b = 8'd64;  #10 
a = 8'd25; b = 8'd65;  #10 
a = 8'd25; b = 8'd66;  #10 
a = 8'd25; b = 8'd67;  #10 
a = 8'd25; b = 8'd68;  #10 
a = 8'd25; b = 8'd69;  #10 
a = 8'd25; b = 8'd70;  #10 
a = 8'd25; b = 8'd71;  #10 
a = 8'd25; b = 8'd72;  #10 
a = 8'd25; b = 8'd73;  #10 
a = 8'd25; b = 8'd74;  #10 
a = 8'd25; b = 8'd75;  #10 
a = 8'd25; b = 8'd76;  #10 
a = 8'd25; b = 8'd77;  #10 
a = 8'd25; b = 8'd78;  #10 
a = 8'd25; b = 8'd79;  #10 
a = 8'd25; b = 8'd80;  #10 
a = 8'd25; b = 8'd81;  #10 
a = 8'd25; b = 8'd82;  #10 
a = 8'd25; b = 8'd83;  #10 
a = 8'd25; b = 8'd84;  #10 
a = 8'd25; b = 8'd85;  #10 
a = 8'd25; b = 8'd86;  #10 
a = 8'd25; b = 8'd87;  #10 
a = 8'd25; b = 8'd88;  #10 
a = 8'd25; b = 8'd89;  #10 
a = 8'd25; b = 8'd90;  #10 
a = 8'd25; b = 8'd91;  #10 
a = 8'd25; b = 8'd92;  #10 
a = 8'd25; b = 8'd93;  #10 
a = 8'd25; b = 8'd94;  #10 
a = 8'd25; b = 8'd95;  #10 
a = 8'd25; b = 8'd96;  #10 
a = 8'd25; b = 8'd97;  #10 
a = 8'd25; b = 8'd98;  #10 
a = 8'd25; b = 8'd99;  #10 
a = 8'd25; b = 8'd100;  #10 
a = 8'd25; b = 8'd101;  #10 
a = 8'd25; b = 8'd102;  #10 
a = 8'd25; b = 8'd103;  #10 
a = 8'd25; b = 8'd104;  #10 
a = 8'd25; b = 8'd105;  #10 
a = 8'd25; b = 8'd106;  #10 
a = 8'd25; b = 8'd107;  #10 
a = 8'd25; b = 8'd108;  #10 
a = 8'd25; b = 8'd109;  #10 
a = 8'd25; b = 8'd110;  #10 
a = 8'd25; b = 8'd111;  #10 
a = 8'd25; b = 8'd112;  #10 
a = 8'd25; b = 8'd113;  #10 
a = 8'd25; b = 8'd114;  #10 
a = 8'd25; b = 8'd115;  #10 
a = 8'd25; b = 8'd116;  #10 
a = 8'd25; b = 8'd117;  #10 
a = 8'd25; b = 8'd118;  #10 
a = 8'd25; b = 8'd119;  #10 
a = 8'd25; b = 8'd120;  #10 
a = 8'd25; b = 8'd121;  #10 
a = 8'd25; b = 8'd122;  #10 
a = 8'd25; b = 8'd123;  #10 
a = 8'd25; b = 8'd124;  #10 
a = 8'd25; b = 8'd125;  #10 
a = 8'd25; b = 8'd126;  #10 
a = 8'd25; b = 8'd127;  #10 
a = 8'd25; b = 8'd128;  #10 
a = 8'd25; b = 8'd129;  #10 
a = 8'd25; b = 8'd130;  #10 
a = 8'd25; b = 8'd131;  #10 
a = 8'd25; b = 8'd132;  #10 
a = 8'd25; b = 8'd133;  #10 
a = 8'd25; b = 8'd134;  #10 
a = 8'd25; b = 8'd135;  #10 
a = 8'd25; b = 8'd136;  #10 
a = 8'd25; b = 8'd137;  #10 
a = 8'd25; b = 8'd138;  #10 
a = 8'd25; b = 8'd139;  #10 
a = 8'd25; b = 8'd140;  #10 
a = 8'd25; b = 8'd141;  #10 
a = 8'd25; b = 8'd142;  #10 
a = 8'd25; b = 8'd143;  #10 
a = 8'd25; b = 8'd144;  #10 
a = 8'd25; b = 8'd145;  #10 
a = 8'd25; b = 8'd146;  #10 
a = 8'd25; b = 8'd147;  #10 
a = 8'd25; b = 8'd148;  #10 
a = 8'd25; b = 8'd149;  #10 
a = 8'd25; b = 8'd150;  #10 
a = 8'd25; b = 8'd151;  #10 
a = 8'd25; b = 8'd152;  #10 
a = 8'd25; b = 8'd153;  #10 
a = 8'd25; b = 8'd154;  #10 
a = 8'd25; b = 8'd155;  #10 
a = 8'd25; b = 8'd156;  #10 
a = 8'd25; b = 8'd157;  #10 
a = 8'd25; b = 8'd158;  #10 
a = 8'd25; b = 8'd159;  #10 
a = 8'd25; b = 8'd160;  #10 
a = 8'd25; b = 8'd161;  #10 
a = 8'd25; b = 8'd162;  #10 
a = 8'd25; b = 8'd163;  #10 
a = 8'd25; b = 8'd164;  #10 
a = 8'd25; b = 8'd165;  #10 
a = 8'd25; b = 8'd166;  #10 
a = 8'd25; b = 8'd167;  #10 
a = 8'd25; b = 8'd168;  #10 
a = 8'd25; b = 8'd169;  #10 
a = 8'd25; b = 8'd170;  #10 
a = 8'd25; b = 8'd171;  #10 
a = 8'd25; b = 8'd172;  #10 
a = 8'd25; b = 8'd173;  #10 
a = 8'd25; b = 8'd174;  #10 
a = 8'd25; b = 8'd175;  #10 
a = 8'd25; b = 8'd176;  #10 
a = 8'd25; b = 8'd177;  #10 
a = 8'd25; b = 8'd178;  #10 
a = 8'd25; b = 8'd179;  #10 
a = 8'd25; b = 8'd180;  #10 
a = 8'd25; b = 8'd181;  #10 
a = 8'd25; b = 8'd182;  #10 
a = 8'd25; b = 8'd183;  #10 
a = 8'd25; b = 8'd184;  #10 
a = 8'd25; b = 8'd185;  #10 
a = 8'd25; b = 8'd186;  #10 
a = 8'd25; b = 8'd187;  #10 
a = 8'd25; b = 8'd188;  #10 
a = 8'd25; b = 8'd189;  #10 
a = 8'd25; b = 8'd190;  #10 
a = 8'd25; b = 8'd191;  #10 
a = 8'd25; b = 8'd192;  #10 
a = 8'd25; b = 8'd193;  #10 
a = 8'd25; b = 8'd194;  #10 
a = 8'd25; b = 8'd195;  #10 
a = 8'd25; b = 8'd196;  #10 
a = 8'd25; b = 8'd197;  #10 
a = 8'd25; b = 8'd198;  #10 
a = 8'd25; b = 8'd199;  #10 
a = 8'd25; b = 8'd200;  #10 
a = 8'd25; b = 8'd201;  #10 
a = 8'd25; b = 8'd202;  #10 
a = 8'd25; b = 8'd203;  #10 
a = 8'd25; b = 8'd204;  #10 
a = 8'd25; b = 8'd205;  #10 
a = 8'd25; b = 8'd206;  #10 
a = 8'd25; b = 8'd207;  #10 
a = 8'd25; b = 8'd208;  #10 
a = 8'd25; b = 8'd209;  #10 
a = 8'd25; b = 8'd210;  #10 
a = 8'd25; b = 8'd211;  #10 
a = 8'd25; b = 8'd212;  #10 
a = 8'd25; b = 8'd213;  #10 
a = 8'd25; b = 8'd214;  #10 
a = 8'd25; b = 8'd215;  #10 
a = 8'd25; b = 8'd216;  #10 
a = 8'd25; b = 8'd217;  #10 
a = 8'd25; b = 8'd218;  #10 
a = 8'd25; b = 8'd219;  #10 
a = 8'd25; b = 8'd220;  #10 
a = 8'd25; b = 8'd221;  #10 
a = 8'd25; b = 8'd222;  #10 
a = 8'd25; b = 8'd223;  #10 
a = 8'd25; b = 8'd224;  #10 
a = 8'd25; b = 8'd225;  #10 
a = 8'd25; b = 8'd226;  #10 
a = 8'd25; b = 8'd227;  #10 
a = 8'd25; b = 8'd228;  #10 
a = 8'd25; b = 8'd229;  #10 
a = 8'd25; b = 8'd230;  #10 
a = 8'd25; b = 8'd231;  #10 
a = 8'd25; b = 8'd232;  #10 
a = 8'd25; b = 8'd233;  #10 
a = 8'd25; b = 8'd234;  #10 
a = 8'd25; b = 8'd235;  #10 
a = 8'd25; b = 8'd236;  #10 
a = 8'd25; b = 8'd237;  #10 
a = 8'd25; b = 8'd238;  #10 
a = 8'd25; b = 8'd239;  #10 
a = 8'd25; b = 8'd240;  #10 
a = 8'd25; b = 8'd241;  #10 
a = 8'd25; b = 8'd242;  #10 
a = 8'd25; b = 8'd243;  #10 
a = 8'd25; b = 8'd244;  #10 
a = 8'd25; b = 8'd245;  #10 
a = 8'd25; b = 8'd246;  #10 
a = 8'd25; b = 8'd247;  #10 
a = 8'd25; b = 8'd248;  #10 
a = 8'd25; b = 8'd249;  #10 
a = 8'd25; b = 8'd250;  #10 
a = 8'd25; b = 8'd251;  #10 
a = 8'd25; b = 8'd252;  #10 
a = 8'd25; b = 8'd253;  #10 
a = 8'd25; b = 8'd254;  #10 
a = 8'd25; b = 8'd255;  #10 
a = 8'd26; b = 8'd0;  #10 
a = 8'd26; b = 8'd1;  #10 
a = 8'd26; b = 8'd2;  #10 
a = 8'd26; b = 8'd3;  #10 
a = 8'd26; b = 8'd4;  #10 
a = 8'd26; b = 8'd5;  #10 
a = 8'd26; b = 8'd6;  #10 
a = 8'd26; b = 8'd7;  #10 
a = 8'd26; b = 8'd8;  #10 
a = 8'd26; b = 8'd9;  #10 
a = 8'd26; b = 8'd10;  #10 
a = 8'd26; b = 8'd11;  #10 
a = 8'd26; b = 8'd12;  #10 
a = 8'd26; b = 8'd13;  #10 
a = 8'd26; b = 8'd14;  #10 
a = 8'd26; b = 8'd15;  #10 
a = 8'd26; b = 8'd16;  #10 
a = 8'd26; b = 8'd17;  #10 
a = 8'd26; b = 8'd18;  #10 
a = 8'd26; b = 8'd19;  #10 
a = 8'd26; b = 8'd20;  #10 
a = 8'd26; b = 8'd21;  #10 
a = 8'd26; b = 8'd22;  #10 
a = 8'd26; b = 8'd23;  #10 
a = 8'd26; b = 8'd24;  #10 
a = 8'd26; b = 8'd25;  #10 
a = 8'd26; b = 8'd26;  #10 
a = 8'd26; b = 8'd27;  #10 
a = 8'd26; b = 8'd28;  #10 
a = 8'd26; b = 8'd29;  #10 
a = 8'd26; b = 8'd30;  #10 
a = 8'd26; b = 8'd31;  #10 
a = 8'd26; b = 8'd32;  #10 
a = 8'd26; b = 8'd33;  #10 
a = 8'd26; b = 8'd34;  #10 
a = 8'd26; b = 8'd35;  #10 
a = 8'd26; b = 8'd36;  #10 
a = 8'd26; b = 8'd37;  #10 
a = 8'd26; b = 8'd38;  #10 
a = 8'd26; b = 8'd39;  #10 
a = 8'd26; b = 8'd40;  #10 
a = 8'd26; b = 8'd41;  #10 
a = 8'd26; b = 8'd42;  #10 
a = 8'd26; b = 8'd43;  #10 
a = 8'd26; b = 8'd44;  #10 
a = 8'd26; b = 8'd45;  #10 
a = 8'd26; b = 8'd46;  #10 
a = 8'd26; b = 8'd47;  #10 
a = 8'd26; b = 8'd48;  #10 
a = 8'd26; b = 8'd49;  #10 
a = 8'd26; b = 8'd50;  #10 
a = 8'd26; b = 8'd51;  #10 
a = 8'd26; b = 8'd52;  #10 
a = 8'd26; b = 8'd53;  #10 
a = 8'd26; b = 8'd54;  #10 
a = 8'd26; b = 8'd55;  #10 
a = 8'd26; b = 8'd56;  #10 
a = 8'd26; b = 8'd57;  #10 
a = 8'd26; b = 8'd58;  #10 
a = 8'd26; b = 8'd59;  #10 
a = 8'd26; b = 8'd60;  #10 
a = 8'd26; b = 8'd61;  #10 
a = 8'd26; b = 8'd62;  #10 
a = 8'd26; b = 8'd63;  #10 
a = 8'd26; b = 8'd64;  #10 
a = 8'd26; b = 8'd65;  #10 
a = 8'd26; b = 8'd66;  #10 
a = 8'd26; b = 8'd67;  #10 
a = 8'd26; b = 8'd68;  #10 
a = 8'd26; b = 8'd69;  #10 
a = 8'd26; b = 8'd70;  #10 
a = 8'd26; b = 8'd71;  #10 
a = 8'd26; b = 8'd72;  #10 
a = 8'd26; b = 8'd73;  #10 
a = 8'd26; b = 8'd74;  #10 
a = 8'd26; b = 8'd75;  #10 
a = 8'd26; b = 8'd76;  #10 
a = 8'd26; b = 8'd77;  #10 
a = 8'd26; b = 8'd78;  #10 
a = 8'd26; b = 8'd79;  #10 
a = 8'd26; b = 8'd80;  #10 
a = 8'd26; b = 8'd81;  #10 
a = 8'd26; b = 8'd82;  #10 
a = 8'd26; b = 8'd83;  #10 
a = 8'd26; b = 8'd84;  #10 
a = 8'd26; b = 8'd85;  #10 
a = 8'd26; b = 8'd86;  #10 
a = 8'd26; b = 8'd87;  #10 
a = 8'd26; b = 8'd88;  #10 
a = 8'd26; b = 8'd89;  #10 
a = 8'd26; b = 8'd90;  #10 
a = 8'd26; b = 8'd91;  #10 
a = 8'd26; b = 8'd92;  #10 
a = 8'd26; b = 8'd93;  #10 
a = 8'd26; b = 8'd94;  #10 
a = 8'd26; b = 8'd95;  #10 
a = 8'd26; b = 8'd96;  #10 
a = 8'd26; b = 8'd97;  #10 
a = 8'd26; b = 8'd98;  #10 
a = 8'd26; b = 8'd99;  #10 
a = 8'd26; b = 8'd100;  #10 
a = 8'd26; b = 8'd101;  #10 
a = 8'd26; b = 8'd102;  #10 
a = 8'd26; b = 8'd103;  #10 
a = 8'd26; b = 8'd104;  #10 
a = 8'd26; b = 8'd105;  #10 
a = 8'd26; b = 8'd106;  #10 
a = 8'd26; b = 8'd107;  #10 
a = 8'd26; b = 8'd108;  #10 
a = 8'd26; b = 8'd109;  #10 
a = 8'd26; b = 8'd110;  #10 
a = 8'd26; b = 8'd111;  #10 
a = 8'd26; b = 8'd112;  #10 
a = 8'd26; b = 8'd113;  #10 
a = 8'd26; b = 8'd114;  #10 
a = 8'd26; b = 8'd115;  #10 
a = 8'd26; b = 8'd116;  #10 
a = 8'd26; b = 8'd117;  #10 
a = 8'd26; b = 8'd118;  #10 
a = 8'd26; b = 8'd119;  #10 
a = 8'd26; b = 8'd120;  #10 
a = 8'd26; b = 8'd121;  #10 
a = 8'd26; b = 8'd122;  #10 
a = 8'd26; b = 8'd123;  #10 
a = 8'd26; b = 8'd124;  #10 
a = 8'd26; b = 8'd125;  #10 
a = 8'd26; b = 8'd126;  #10 
a = 8'd26; b = 8'd127;  #10 
a = 8'd26; b = 8'd128;  #10 
a = 8'd26; b = 8'd129;  #10 
a = 8'd26; b = 8'd130;  #10 
a = 8'd26; b = 8'd131;  #10 
a = 8'd26; b = 8'd132;  #10 
a = 8'd26; b = 8'd133;  #10 
a = 8'd26; b = 8'd134;  #10 
a = 8'd26; b = 8'd135;  #10 
a = 8'd26; b = 8'd136;  #10 
a = 8'd26; b = 8'd137;  #10 
a = 8'd26; b = 8'd138;  #10 
a = 8'd26; b = 8'd139;  #10 
a = 8'd26; b = 8'd140;  #10 
a = 8'd26; b = 8'd141;  #10 
a = 8'd26; b = 8'd142;  #10 
a = 8'd26; b = 8'd143;  #10 
a = 8'd26; b = 8'd144;  #10 
a = 8'd26; b = 8'd145;  #10 
a = 8'd26; b = 8'd146;  #10 
a = 8'd26; b = 8'd147;  #10 
a = 8'd26; b = 8'd148;  #10 
a = 8'd26; b = 8'd149;  #10 
a = 8'd26; b = 8'd150;  #10 
a = 8'd26; b = 8'd151;  #10 
a = 8'd26; b = 8'd152;  #10 
a = 8'd26; b = 8'd153;  #10 
a = 8'd26; b = 8'd154;  #10 
a = 8'd26; b = 8'd155;  #10 
a = 8'd26; b = 8'd156;  #10 
a = 8'd26; b = 8'd157;  #10 
a = 8'd26; b = 8'd158;  #10 
a = 8'd26; b = 8'd159;  #10 
a = 8'd26; b = 8'd160;  #10 
a = 8'd26; b = 8'd161;  #10 
a = 8'd26; b = 8'd162;  #10 
a = 8'd26; b = 8'd163;  #10 
a = 8'd26; b = 8'd164;  #10 
a = 8'd26; b = 8'd165;  #10 
a = 8'd26; b = 8'd166;  #10 
a = 8'd26; b = 8'd167;  #10 
a = 8'd26; b = 8'd168;  #10 
a = 8'd26; b = 8'd169;  #10 
a = 8'd26; b = 8'd170;  #10 
a = 8'd26; b = 8'd171;  #10 
a = 8'd26; b = 8'd172;  #10 
a = 8'd26; b = 8'd173;  #10 
a = 8'd26; b = 8'd174;  #10 
a = 8'd26; b = 8'd175;  #10 
a = 8'd26; b = 8'd176;  #10 
a = 8'd26; b = 8'd177;  #10 
a = 8'd26; b = 8'd178;  #10 
a = 8'd26; b = 8'd179;  #10 
a = 8'd26; b = 8'd180;  #10 
a = 8'd26; b = 8'd181;  #10 
a = 8'd26; b = 8'd182;  #10 
a = 8'd26; b = 8'd183;  #10 
a = 8'd26; b = 8'd184;  #10 
a = 8'd26; b = 8'd185;  #10 
a = 8'd26; b = 8'd186;  #10 
a = 8'd26; b = 8'd187;  #10 
a = 8'd26; b = 8'd188;  #10 
a = 8'd26; b = 8'd189;  #10 
a = 8'd26; b = 8'd190;  #10 
a = 8'd26; b = 8'd191;  #10 
a = 8'd26; b = 8'd192;  #10 
a = 8'd26; b = 8'd193;  #10 
a = 8'd26; b = 8'd194;  #10 
a = 8'd26; b = 8'd195;  #10 
a = 8'd26; b = 8'd196;  #10 
a = 8'd26; b = 8'd197;  #10 
a = 8'd26; b = 8'd198;  #10 
a = 8'd26; b = 8'd199;  #10 
a = 8'd26; b = 8'd200;  #10 
a = 8'd26; b = 8'd201;  #10 
a = 8'd26; b = 8'd202;  #10 
a = 8'd26; b = 8'd203;  #10 
a = 8'd26; b = 8'd204;  #10 
a = 8'd26; b = 8'd205;  #10 
a = 8'd26; b = 8'd206;  #10 
a = 8'd26; b = 8'd207;  #10 
a = 8'd26; b = 8'd208;  #10 
a = 8'd26; b = 8'd209;  #10 
a = 8'd26; b = 8'd210;  #10 
a = 8'd26; b = 8'd211;  #10 
a = 8'd26; b = 8'd212;  #10 
a = 8'd26; b = 8'd213;  #10 
a = 8'd26; b = 8'd214;  #10 
a = 8'd26; b = 8'd215;  #10 
a = 8'd26; b = 8'd216;  #10 
a = 8'd26; b = 8'd217;  #10 
a = 8'd26; b = 8'd218;  #10 
a = 8'd26; b = 8'd219;  #10 
a = 8'd26; b = 8'd220;  #10 
a = 8'd26; b = 8'd221;  #10 
a = 8'd26; b = 8'd222;  #10 
a = 8'd26; b = 8'd223;  #10 
a = 8'd26; b = 8'd224;  #10 
a = 8'd26; b = 8'd225;  #10 
a = 8'd26; b = 8'd226;  #10 
a = 8'd26; b = 8'd227;  #10 
a = 8'd26; b = 8'd228;  #10 
a = 8'd26; b = 8'd229;  #10 
a = 8'd26; b = 8'd230;  #10 
a = 8'd26; b = 8'd231;  #10 
a = 8'd26; b = 8'd232;  #10 
a = 8'd26; b = 8'd233;  #10 
a = 8'd26; b = 8'd234;  #10 
a = 8'd26; b = 8'd235;  #10 
a = 8'd26; b = 8'd236;  #10 
a = 8'd26; b = 8'd237;  #10 
a = 8'd26; b = 8'd238;  #10 
a = 8'd26; b = 8'd239;  #10 
a = 8'd26; b = 8'd240;  #10 
a = 8'd26; b = 8'd241;  #10 
a = 8'd26; b = 8'd242;  #10 
a = 8'd26; b = 8'd243;  #10 
a = 8'd26; b = 8'd244;  #10 
a = 8'd26; b = 8'd245;  #10 
a = 8'd26; b = 8'd246;  #10 
a = 8'd26; b = 8'd247;  #10 
a = 8'd26; b = 8'd248;  #10 
a = 8'd26; b = 8'd249;  #10 
a = 8'd26; b = 8'd250;  #10 
a = 8'd26; b = 8'd251;  #10 
a = 8'd26; b = 8'd252;  #10 
a = 8'd26; b = 8'd253;  #10 
a = 8'd26; b = 8'd254;  #10 
a = 8'd26; b = 8'd255;  #10 
a = 8'd27; b = 8'd0;  #10 
a = 8'd27; b = 8'd1;  #10 
a = 8'd27; b = 8'd2;  #10 
a = 8'd27; b = 8'd3;  #10 
a = 8'd27; b = 8'd4;  #10 
a = 8'd27; b = 8'd5;  #10 
a = 8'd27; b = 8'd6;  #10 
a = 8'd27; b = 8'd7;  #10 
a = 8'd27; b = 8'd8;  #10 
a = 8'd27; b = 8'd9;  #10 
a = 8'd27; b = 8'd10;  #10 
a = 8'd27; b = 8'd11;  #10 
a = 8'd27; b = 8'd12;  #10 
a = 8'd27; b = 8'd13;  #10 
a = 8'd27; b = 8'd14;  #10 
a = 8'd27; b = 8'd15;  #10 
a = 8'd27; b = 8'd16;  #10 
a = 8'd27; b = 8'd17;  #10 
a = 8'd27; b = 8'd18;  #10 
a = 8'd27; b = 8'd19;  #10 
a = 8'd27; b = 8'd20;  #10 
a = 8'd27; b = 8'd21;  #10 
a = 8'd27; b = 8'd22;  #10 
a = 8'd27; b = 8'd23;  #10 
a = 8'd27; b = 8'd24;  #10 
a = 8'd27; b = 8'd25;  #10 
a = 8'd27; b = 8'd26;  #10 
a = 8'd27; b = 8'd27;  #10 
a = 8'd27; b = 8'd28;  #10 
a = 8'd27; b = 8'd29;  #10 
a = 8'd27; b = 8'd30;  #10 
a = 8'd27; b = 8'd31;  #10 
a = 8'd27; b = 8'd32;  #10 
a = 8'd27; b = 8'd33;  #10 
a = 8'd27; b = 8'd34;  #10 
a = 8'd27; b = 8'd35;  #10 
a = 8'd27; b = 8'd36;  #10 
a = 8'd27; b = 8'd37;  #10 
a = 8'd27; b = 8'd38;  #10 
a = 8'd27; b = 8'd39;  #10 
a = 8'd27; b = 8'd40;  #10 
a = 8'd27; b = 8'd41;  #10 
a = 8'd27; b = 8'd42;  #10 
a = 8'd27; b = 8'd43;  #10 
a = 8'd27; b = 8'd44;  #10 
a = 8'd27; b = 8'd45;  #10 
a = 8'd27; b = 8'd46;  #10 
a = 8'd27; b = 8'd47;  #10 
a = 8'd27; b = 8'd48;  #10 
a = 8'd27; b = 8'd49;  #10 
a = 8'd27; b = 8'd50;  #10 
a = 8'd27; b = 8'd51;  #10 
a = 8'd27; b = 8'd52;  #10 
a = 8'd27; b = 8'd53;  #10 
a = 8'd27; b = 8'd54;  #10 
a = 8'd27; b = 8'd55;  #10 
a = 8'd27; b = 8'd56;  #10 
a = 8'd27; b = 8'd57;  #10 
a = 8'd27; b = 8'd58;  #10 
a = 8'd27; b = 8'd59;  #10 
a = 8'd27; b = 8'd60;  #10 
a = 8'd27; b = 8'd61;  #10 
a = 8'd27; b = 8'd62;  #10 
a = 8'd27; b = 8'd63;  #10 
a = 8'd27; b = 8'd64;  #10 
a = 8'd27; b = 8'd65;  #10 
a = 8'd27; b = 8'd66;  #10 
a = 8'd27; b = 8'd67;  #10 
a = 8'd27; b = 8'd68;  #10 
a = 8'd27; b = 8'd69;  #10 
a = 8'd27; b = 8'd70;  #10 
a = 8'd27; b = 8'd71;  #10 
a = 8'd27; b = 8'd72;  #10 
a = 8'd27; b = 8'd73;  #10 
a = 8'd27; b = 8'd74;  #10 
a = 8'd27; b = 8'd75;  #10 
a = 8'd27; b = 8'd76;  #10 
a = 8'd27; b = 8'd77;  #10 
a = 8'd27; b = 8'd78;  #10 
a = 8'd27; b = 8'd79;  #10 
a = 8'd27; b = 8'd80;  #10 
a = 8'd27; b = 8'd81;  #10 
a = 8'd27; b = 8'd82;  #10 
a = 8'd27; b = 8'd83;  #10 
a = 8'd27; b = 8'd84;  #10 
a = 8'd27; b = 8'd85;  #10 
a = 8'd27; b = 8'd86;  #10 
a = 8'd27; b = 8'd87;  #10 
a = 8'd27; b = 8'd88;  #10 
a = 8'd27; b = 8'd89;  #10 
a = 8'd27; b = 8'd90;  #10 
a = 8'd27; b = 8'd91;  #10 
a = 8'd27; b = 8'd92;  #10 
a = 8'd27; b = 8'd93;  #10 
a = 8'd27; b = 8'd94;  #10 
a = 8'd27; b = 8'd95;  #10 
a = 8'd27; b = 8'd96;  #10 
a = 8'd27; b = 8'd97;  #10 
a = 8'd27; b = 8'd98;  #10 
a = 8'd27; b = 8'd99;  #10 
a = 8'd27; b = 8'd100;  #10 
a = 8'd27; b = 8'd101;  #10 
a = 8'd27; b = 8'd102;  #10 
a = 8'd27; b = 8'd103;  #10 
a = 8'd27; b = 8'd104;  #10 
a = 8'd27; b = 8'd105;  #10 
a = 8'd27; b = 8'd106;  #10 
a = 8'd27; b = 8'd107;  #10 
a = 8'd27; b = 8'd108;  #10 
a = 8'd27; b = 8'd109;  #10 
a = 8'd27; b = 8'd110;  #10 
a = 8'd27; b = 8'd111;  #10 
a = 8'd27; b = 8'd112;  #10 
a = 8'd27; b = 8'd113;  #10 
a = 8'd27; b = 8'd114;  #10 
a = 8'd27; b = 8'd115;  #10 
a = 8'd27; b = 8'd116;  #10 
a = 8'd27; b = 8'd117;  #10 
a = 8'd27; b = 8'd118;  #10 
a = 8'd27; b = 8'd119;  #10 
a = 8'd27; b = 8'd120;  #10 
a = 8'd27; b = 8'd121;  #10 
a = 8'd27; b = 8'd122;  #10 
a = 8'd27; b = 8'd123;  #10 
a = 8'd27; b = 8'd124;  #10 
a = 8'd27; b = 8'd125;  #10 
a = 8'd27; b = 8'd126;  #10 
a = 8'd27; b = 8'd127;  #10 
a = 8'd27; b = 8'd128;  #10 
a = 8'd27; b = 8'd129;  #10 
a = 8'd27; b = 8'd130;  #10 
a = 8'd27; b = 8'd131;  #10 
a = 8'd27; b = 8'd132;  #10 
a = 8'd27; b = 8'd133;  #10 
a = 8'd27; b = 8'd134;  #10 
a = 8'd27; b = 8'd135;  #10 
a = 8'd27; b = 8'd136;  #10 
a = 8'd27; b = 8'd137;  #10 
a = 8'd27; b = 8'd138;  #10 
a = 8'd27; b = 8'd139;  #10 
a = 8'd27; b = 8'd140;  #10 
a = 8'd27; b = 8'd141;  #10 
a = 8'd27; b = 8'd142;  #10 
a = 8'd27; b = 8'd143;  #10 
a = 8'd27; b = 8'd144;  #10 
a = 8'd27; b = 8'd145;  #10 
a = 8'd27; b = 8'd146;  #10 
a = 8'd27; b = 8'd147;  #10 
a = 8'd27; b = 8'd148;  #10 
a = 8'd27; b = 8'd149;  #10 
a = 8'd27; b = 8'd150;  #10 
a = 8'd27; b = 8'd151;  #10 
a = 8'd27; b = 8'd152;  #10 
a = 8'd27; b = 8'd153;  #10 
a = 8'd27; b = 8'd154;  #10 
a = 8'd27; b = 8'd155;  #10 
a = 8'd27; b = 8'd156;  #10 
a = 8'd27; b = 8'd157;  #10 
a = 8'd27; b = 8'd158;  #10 
a = 8'd27; b = 8'd159;  #10 
a = 8'd27; b = 8'd160;  #10 
a = 8'd27; b = 8'd161;  #10 
a = 8'd27; b = 8'd162;  #10 
a = 8'd27; b = 8'd163;  #10 
a = 8'd27; b = 8'd164;  #10 
a = 8'd27; b = 8'd165;  #10 
a = 8'd27; b = 8'd166;  #10 
a = 8'd27; b = 8'd167;  #10 
a = 8'd27; b = 8'd168;  #10 
a = 8'd27; b = 8'd169;  #10 
a = 8'd27; b = 8'd170;  #10 
a = 8'd27; b = 8'd171;  #10 
a = 8'd27; b = 8'd172;  #10 
a = 8'd27; b = 8'd173;  #10 
a = 8'd27; b = 8'd174;  #10 
a = 8'd27; b = 8'd175;  #10 
a = 8'd27; b = 8'd176;  #10 
a = 8'd27; b = 8'd177;  #10 
a = 8'd27; b = 8'd178;  #10 
a = 8'd27; b = 8'd179;  #10 
a = 8'd27; b = 8'd180;  #10 
a = 8'd27; b = 8'd181;  #10 
a = 8'd27; b = 8'd182;  #10 
a = 8'd27; b = 8'd183;  #10 
a = 8'd27; b = 8'd184;  #10 
a = 8'd27; b = 8'd185;  #10 
a = 8'd27; b = 8'd186;  #10 
a = 8'd27; b = 8'd187;  #10 
a = 8'd27; b = 8'd188;  #10 
a = 8'd27; b = 8'd189;  #10 
a = 8'd27; b = 8'd190;  #10 
a = 8'd27; b = 8'd191;  #10 
a = 8'd27; b = 8'd192;  #10 
a = 8'd27; b = 8'd193;  #10 
a = 8'd27; b = 8'd194;  #10 
a = 8'd27; b = 8'd195;  #10 
a = 8'd27; b = 8'd196;  #10 
a = 8'd27; b = 8'd197;  #10 
a = 8'd27; b = 8'd198;  #10 
a = 8'd27; b = 8'd199;  #10 
a = 8'd27; b = 8'd200;  #10 
a = 8'd27; b = 8'd201;  #10 
a = 8'd27; b = 8'd202;  #10 
a = 8'd27; b = 8'd203;  #10 
a = 8'd27; b = 8'd204;  #10 
a = 8'd27; b = 8'd205;  #10 
a = 8'd27; b = 8'd206;  #10 
a = 8'd27; b = 8'd207;  #10 
a = 8'd27; b = 8'd208;  #10 
a = 8'd27; b = 8'd209;  #10 
a = 8'd27; b = 8'd210;  #10 
a = 8'd27; b = 8'd211;  #10 
a = 8'd27; b = 8'd212;  #10 
a = 8'd27; b = 8'd213;  #10 
a = 8'd27; b = 8'd214;  #10 
a = 8'd27; b = 8'd215;  #10 
a = 8'd27; b = 8'd216;  #10 
a = 8'd27; b = 8'd217;  #10 
a = 8'd27; b = 8'd218;  #10 
a = 8'd27; b = 8'd219;  #10 
a = 8'd27; b = 8'd220;  #10 
a = 8'd27; b = 8'd221;  #10 
a = 8'd27; b = 8'd222;  #10 
a = 8'd27; b = 8'd223;  #10 
a = 8'd27; b = 8'd224;  #10 
a = 8'd27; b = 8'd225;  #10 
a = 8'd27; b = 8'd226;  #10 
a = 8'd27; b = 8'd227;  #10 
a = 8'd27; b = 8'd228;  #10 
a = 8'd27; b = 8'd229;  #10 
a = 8'd27; b = 8'd230;  #10 
a = 8'd27; b = 8'd231;  #10 
a = 8'd27; b = 8'd232;  #10 
a = 8'd27; b = 8'd233;  #10 
a = 8'd27; b = 8'd234;  #10 
a = 8'd27; b = 8'd235;  #10 
a = 8'd27; b = 8'd236;  #10 
a = 8'd27; b = 8'd237;  #10 
a = 8'd27; b = 8'd238;  #10 
a = 8'd27; b = 8'd239;  #10 
a = 8'd27; b = 8'd240;  #10 
a = 8'd27; b = 8'd241;  #10 
a = 8'd27; b = 8'd242;  #10 
a = 8'd27; b = 8'd243;  #10 
a = 8'd27; b = 8'd244;  #10 
a = 8'd27; b = 8'd245;  #10 
a = 8'd27; b = 8'd246;  #10 
a = 8'd27; b = 8'd247;  #10 
a = 8'd27; b = 8'd248;  #10 
a = 8'd27; b = 8'd249;  #10 
a = 8'd27; b = 8'd250;  #10 
a = 8'd27; b = 8'd251;  #10 
a = 8'd27; b = 8'd252;  #10 
a = 8'd27; b = 8'd253;  #10 
a = 8'd27; b = 8'd254;  #10 
a = 8'd27; b = 8'd255;  #10 
a = 8'd28; b = 8'd0;  #10 
a = 8'd28; b = 8'd1;  #10 
a = 8'd28; b = 8'd2;  #10 
a = 8'd28; b = 8'd3;  #10 
a = 8'd28; b = 8'd4;  #10 
a = 8'd28; b = 8'd5;  #10 
a = 8'd28; b = 8'd6;  #10 
a = 8'd28; b = 8'd7;  #10 
a = 8'd28; b = 8'd8;  #10 
a = 8'd28; b = 8'd9;  #10 
a = 8'd28; b = 8'd10;  #10 
a = 8'd28; b = 8'd11;  #10 
a = 8'd28; b = 8'd12;  #10 
a = 8'd28; b = 8'd13;  #10 
a = 8'd28; b = 8'd14;  #10 
a = 8'd28; b = 8'd15;  #10 
a = 8'd28; b = 8'd16;  #10 
a = 8'd28; b = 8'd17;  #10 
a = 8'd28; b = 8'd18;  #10 
a = 8'd28; b = 8'd19;  #10 
a = 8'd28; b = 8'd20;  #10 
a = 8'd28; b = 8'd21;  #10 
a = 8'd28; b = 8'd22;  #10 
a = 8'd28; b = 8'd23;  #10 
a = 8'd28; b = 8'd24;  #10 
a = 8'd28; b = 8'd25;  #10 
a = 8'd28; b = 8'd26;  #10 
a = 8'd28; b = 8'd27;  #10 
a = 8'd28; b = 8'd28;  #10 
a = 8'd28; b = 8'd29;  #10 
a = 8'd28; b = 8'd30;  #10 
a = 8'd28; b = 8'd31;  #10 
a = 8'd28; b = 8'd32;  #10 
a = 8'd28; b = 8'd33;  #10 
a = 8'd28; b = 8'd34;  #10 
a = 8'd28; b = 8'd35;  #10 
a = 8'd28; b = 8'd36;  #10 
a = 8'd28; b = 8'd37;  #10 
a = 8'd28; b = 8'd38;  #10 
a = 8'd28; b = 8'd39;  #10 
a = 8'd28; b = 8'd40;  #10 
a = 8'd28; b = 8'd41;  #10 
a = 8'd28; b = 8'd42;  #10 
a = 8'd28; b = 8'd43;  #10 
a = 8'd28; b = 8'd44;  #10 
a = 8'd28; b = 8'd45;  #10 
a = 8'd28; b = 8'd46;  #10 
a = 8'd28; b = 8'd47;  #10 
a = 8'd28; b = 8'd48;  #10 
a = 8'd28; b = 8'd49;  #10 
a = 8'd28; b = 8'd50;  #10 
a = 8'd28; b = 8'd51;  #10 
a = 8'd28; b = 8'd52;  #10 
a = 8'd28; b = 8'd53;  #10 
a = 8'd28; b = 8'd54;  #10 
a = 8'd28; b = 8'd55;  #10 
a = 8'd28; b = 8'd56;  #10 
a = 8'd28; b = 8'd57;  #10 
a = 8'd28; b = 8'd58;  #10 
a = 8'd28; b = 8'd59;  #10 
a = 8'd28; b = 8'd60;  #10 
a = 8'd28; b = 8'd61;  #10 
a = 8'd28; b = 8'd62;  #10 
a = 8'd28; b = 8'd63;  #10 
a = 8'd28; b = 8'd64;  #10 
a = 8'd28; b = 8'd65;  #10 
a = 8'd28; b = 8'd66;  #10 
a = 8'd28; b = 8'd67;  #10 
a = 8'd28; b = 8'd68;  #10 
a = 8'd28; b = 8'd69;  #10 
a = 8'd28; b = 8'd70;  #10 
a = 8'd28; b = 8'd71;  #10 
a = 8'd28; b = 8'd72;  #10 
a = 8'd28; b = 8'd73;  #10 
a = 8'd28; b = 8'd74;  #10 
a = 8'd28; b = 8'd75;  #10 
a = 8'd28; b = 8'd76;  #10 
a = 8'd28; b = 8'd77;  #10 
a = 8'd28; b = 8'd78;  #10 
a = 8'd28; b = 8'd79;  #10 
a = 8'd28; b = 8'd80;  #10 
a = 8'd28; b = 8'd81;  #10 
a = 8'd28; b = 8'd82;  #10 
a = 8'd28; b = 8'd83;  #10 
a = 8'd28; b = 8'd84;  #10 
a = 8'd28; b = 8'd85;  #10 
a = 8'd28; b = 8'd86;  #10 
a = 8'd28; b = 8'd87;  #10 
a = 8'd28; b = 8'd88;  #10 
a = 8'd28; b = 8'd89;  #10 
a = 8'd28; b = 8'd90;  #10 
a = 8'd28; b = 8'd91;  #10 
a = 8'd28; b = 8'd92;  #10 
a = 8'd28; b = 8'd93;  #10 
a = 8'd28; b = 8'd94;  #10 
a = 8'd28; b = 8'd95;  #10 
a = 8'd28; b = 8'd96;  #10 
a = 8'd28; b = 8'd97;  #10 
a = 8'd28; b = 8'd98;  #10 
a = 8'd28; b = 8'd99;  #10 
a = 8'd28; b = 8'd100;  #10 
a = 8'd28; b = 8'd101;  #10 
a = 8'd28; b = 8'd102;  #10 
a = 8'd28; b = 8'd103;  #10 
a = 8'd28; b = 8'd104;  #10 
a = 8'd28; b = 8'd105;  #10 
a = 8'd28; b = 8'd106;  #10 
a = 8'd28; b = 8'd107;  #10 
a = 8'd28; b = 8'd108;  #10 
a = 8'd28; b = 8'd109;  #10 
a = 8'd28; b = 8'd110;  #10 
a = 8'd28; b = 8'd111;  #10 
a = 8'd28; b = 8'd112;  #10 
a = 8'd28; b = 8'd113;  #10 
a = 8'd28; b = 8'd114;  #10 
a = 8'd28; b = 8'd115;  #10 
a = 8'd28; b = 8'd116;  #10 
a = 8'd28; b = 8'd117;  #10 
a = 8'd28; b = 8'd118;  #10 
a = 8'd28; b = 8'd119;  #10 
a = 8'd28; b = 8'd120;  #10 
a = 8'd28; b = 8'd121;  #10 
a = 8'd28; b = 8'd122;  #10 
a = 8'd28; b = 8'd123;  #10 
a = 8'd28; b = 8'd124;  #10 
a = 8'd28; b = 8'd125;  #10 
a = 8'd28; b = 8'd126;  #10 
a = 8'd28; b = 8'd127;  #10 
a = 8'd28; b = 8'd128;  #10 
a = 8'd28; b = 8'd129;  #10 
a = 8'd28; b = 8'd130;  #10 
a = 8'd28; b = 8'd131;  #10 
a = 8'd28; b = 8'd132;  #10 
a = 8'd28; b = 8'd133;  #10 
a = 8'd28; b = 8'd134;  #10 
a = 8'd28; b = 8'd135;  #10 
a = 8'd28; b = 8'd136;  #10 
a = 8'd28; b = 8'd137;  #10 
a = 8'd28; b = 8'd138;  #10 
a = 8'd28; b = 8'd139;  #10 
a = 8'd28; b = 8'd140;  #10 
a = 8'd28; b = 8'd141;  #10 
a = 8'd28; b = 8'd142;  #10 
a = 8'd28; b = 8'd143;  #10 
a = 8'd28; b = 8'd144;  #10 
a = 8'd28; b = 8'd145;  #10 
a = 8'd28; b = 8'd146;  #10 
a = 8'd28; b = 8'd147;  #10 
a = 8'd28; b = 8'd148;  #10 
a = 8'd28; b = 8'd149;  #10 
a = 8'd28; b = 8'd150;  #10 
a = 8'd28; b = 8'd151;  #10 
a = 8'd28; b = 8'd152;  #10 
a = 8'd28; b = 8'd153;  #10 
a = 8'd28; b = 8'd154;  #10 
a = 8'd28; b = 8'd155;  #10 
a = 8'd28; b = 8'd156;  #10 
a = 8'd28; b = 8'd157;  #10 
a = 8'd28; b = 8'd158;  #10 
a = 8'd28; b = 8'd159;  #10 
a = 8'd28; b = 8'd160;  #10 
a = 8'd28; b = 8'd161;  #10 
a = 8'd28; b = 8'd162;  #10 
a = 8'd28; b = 8'd163;  #10 
a = 8'd28; b = 8'd164;  #10 
a = 8'd28; b = 8'd165;  #10 
a = 8'd28; b = 8'd166;  #10 
a = 8'd28; b = 8'd167;  #10 
a = 8'd28; b = 8'd168;  #10 
a = 8'd28; b = 8'd169;  #10 
a = 8'd28; b = 8'd170;  #10 
a = 8'd28; b = 8'd171;  #10 
a = 8'd28; b = 8'd172;  #10 
a = 8'd28; b = 8'd173;  #10 
a = 8'd28; b = 8'd174;  #10 
a = 8'd28; b = 8'd175;  #10 
a = 8'd28; b = 8'd176;  #10 
a = 8'd28; b = 8'd177;  #10 
a = 8'd28; b = 8'd178;  #10 
a = 8'd28; b = 8'd179;  #10 
a = 8'd28; b = 8'd180;  #10 
a = 8'd28; b = 8'd181;  #10 
a = 8'd28; b = 8'd182;  #10 
a = 8'd28; b = 8'd183;  #10 
a = 8'd28; b = 8'd184;  #10 
a = 8'd28; b = 8'd185;  #10 
a = 8'd28; b = 8'd186;  #10 
a = 8'd28; b = 8'd187;  #10 
a = 8'd28; b = 8'd188;  #10 
a = 8'd28; b = 8'd189;  #10 
a = 8'd28; b = 8'd190;  #10 
a = 8'd28; b = 8'd191;  #10 
a = 8'd28; b = 8'd192;  #10 
a = 8'd28; b = 8'd193;  #10 
a = 8'd28; b = 8'd194;  #10 
a = 8'd28; b = 8'd195;  #10 
a = 8'd28; b = 8'd196;  #10 
a = 8'd28; b = 8'd197;  #10 
a = 8'd28; b = 8'd198;  #10 
a = 8'd28; b = 8'd199;  #10 
a = 8'd28; b = 8'd200;  #10 
a = 8'd28; b = 8'd201;  #10 
a = 8'd28; b = 8'd202;  #10 
a = 8'd28; b = 8'd203;  #10 
a = 8'd28; b = 8'd204;  #10 
a = 8'd28; b = 8'd205;  #10 
a = 8'd28; b = 8'd206;  #10 
a = 8'd28; b = 8'd207;  #10 
a = 8'd28; b = 8'd208;  #10 
a = 8'd28; b = 8'd209;  #10 
a = 8'd28; b = 8'd210;  #10 
a = 8'd28; b = 8'd211;  #10 
a = 8'd28; b = 8'd212;  #10 
a = 8'd28; b = 8'd213;  #10 
a = 8'd28; b = 8'd214;  #10 
a = 8'd28; b = 8'd215;  #10 
a = 8'd28; b = 8'd216;  #10 
a = 8'd28; b = 8'd217;  #10 
a = 8'd28; b = 8'd218;  #10 
a = 8'd28; b = 8'd219;  #10 
a = 8'd28; b = 8'd220;  #10 
a = 8'd28; b = 8'd221;  #10 
a = 8'd28; b = 8'd222;  #10 
a = 8'd28; b = 8'd223;  #10 
a = 8'd28; b = 8'd224;  #10 
a = 8'd28; b = 8'd225;  #10 
a = 8'd28; b = 8'd226;  #10 
a = 8'd28; b = 8'd227;  #10 
a = 8'd28; b = 8'd228;  #10 
a = 8'd28; b = 8'd229;  #10 
a = 8'd28; b = 8'd230;  #10 
a = 8'd28; b = 8'd231;  #10 
a = 8'd28; b = 8'd232;  #10 
a = 8'd28; b = 8'd233;  #10 
a = 8'd28; b = 8'd234;  #10 
a = 8'd28; b = 8'd235;  #10 
a = 8'd28; b = 8'd236;  #10 
a = 8'd28; b = 8'd237;  #10 
a = 8'd28; b = 8'd238;  #10 
a = 8'd28; b = 8'd239;  #10 
a = 8'd28; b = 8'd240;  #10 
a = 8'd28; b = 8'd241;  #10 
a = 8'd28; b = 8'd242;  #10 
a = 8'd28; b = 8'd243;  #10 
a = 8'd28; b = 8'd244;  #10 
a = 8'd28; b = 8'd245;  #10 
a = 8'd28; b = 8'd246;  #10 
a = 8'd28; b = 8'd247;  #10 
a = 8'd28; b = 8'd248;  #10 
a = 8'd28; b = 8'd249;  #10 
a = 8'd28; b = 8'd250;  #10 
a = 8'd28; b = 8'd251;  #10 
a = 8'd28; b = 8'd252;  #10 
a = 8'd28; b = 8'd253;  #10 
a = 8'd28; b = 8'd254;  #10 
a = 8'd28; b = 8'd255;  #10 
a = 8'd29; b = 8'd0;  #10 
a = 8'd29; b = 8'd1;  #10 
a = 8'd29; b = 8'd2;  #10 
a = 8'd29; b = 8'd3;  #10 
a = 8'd29; b = 8'd4;  #10 
a = 8'd29; b = 8'd5;  #10 
a = 8'd29; b = 8'd6;  #10 
a = 8'd29; b = 8'd7;  #10 
a = 8'd29; b = 8'd8;  #10 
a = 8'd29; b = 8'd9;  #10 
a = 8'd29; b = 8'd10;  #10 
a = 8'd29; b = 8'd11;  #10 
a = 8'd29; b = 8'd12;  #10 
a = 8'd29; b = 8'd13;  #10 
a = 8'd29; b = 8'd14;  #10 
a = 8'd29; b = 8'd15;  #10 
a = 8'd29; b = 8'd16;  #10 
a = 8'd29; b = 8'd17;  #10 
a = 8'd29; b = 8'd18;  #10 
a = 8'd29; b = 8'd19;  #10 
a = 8'd29; b = 8'd20;  #10 
a = 8'd29; b = 8'd21;  #10 
a = 8'd29; b = 8'd22;  #10 
a = 8'd29; b = 8'd23;  #10 
a = 8'd29; b = 8'd24;  #10 
a = 8'd29; b = 8'd25;  #10 
a = 8'd29; b = 8'd26;  #10 
a = 8'd29; b = 8'd27;  #10 
a = 8'd29; b = 8'd28;  #10 
a = 8'd29; b = 8'd29;  #10 
a = 8'd29; b = 8'd30;  #10 
a = 8'd29; b = 8'd31;  #10 
a = 8'd29; b = 8'd32;  #10 
a = 8'd29; b = 8'd33;  #10 
a = 8'd29; b = 8'd34;  #10 
a = 8'd29; b = 8'd35;  #10 
a = 8'd29; b = 8'd36;  #10 
a = 8'd29; b = 8'd37;  #10 
a = 8'd29; b = 8'd38;  #10 
a = 8'd29; b = 8'd39;  #10 
a = 8'd29; b = 8'd40;  #10 
a = 8'd29; b = 8'd41;  #10 
a = 8'd29; b = 8'd42;  #10 
a = 8'd29; b = 8'd43;  #10 
a = 8'd29; b = 8'd44;  #10 
a = 8'd29; b = 8'd45;  #10 
a = 8'd29; b = 8'd46;  #10 
a = 8'd29; b = 8'd47;  #10 
a = 8'd29; b = 8'd48;  #10 
a = 8'd29; b = 8'd49;  #10 
a = 8'd29; b = 8'd50;  #10 
a = 8'd29; b = 8'd51;  #10 
a = 8'd29; b = 8'd52;  #10 
a = 8'd29; b = 8'd53;  #10 
a = 8'd29; b = 8'd54;  #10 
a = 8'd29; b = 8'd55;  #10 
a = 8'd29; b = 8'd56;  #10 
a = 8'd29; b = 8'd57;  #10 
a = 8'd29; b = 8'd58;  #10 
a = 8'd29; b = 8'd59;  #10 
a = 8'd29; b = 8'd60;  #10 
a = 8'd29; b = 8'd61;  #10 
a = 8'd29; b = 8'd62;  #10 
a = 8'd29; b = 8'd63;  #10 
a = 8'd29; b = 8'd64;  #10 
a = 8'd29; b = 8'd65;  #10 
a = 8'd29; b = 8'd66;  #10 
a = 8'd29; b = 8'd67;  #10 
a = 8'd29; b = 8'd68;  #10 
a = 8'd29; b = 8'd69;  #10 
a = 8'd29; b = 8'd70;  #10 
a = 8'd29; b = 8'd71;  #10 
a = 8'd29; b = 8'd72;  #10 
a = 8'd29; b = 8'd73;  #10 
a = 8'd29; b = 8'd74;  #10 
a = 8'd29; b = 8'd75;  #10 
a = 8'd29; b = 8'd76;  #10 
a = 8'd29; b = 8'd77;  #10 
a = 8'd29; b = 8'd78;  #10 
a = 8'd29; b = 8'd79;  #10 
a = 8'd29; b = 8'd80;  #10 
a = 8'd29; b = 8'd81;  #10 
a = 8'd29; b = 8'd82;  #10 
a = 8'd29; b = 8'd83;  #10 
a = 8'd29; b = 8'd84;  #10 
a = 8'd29; b = 8'd85;  #10 
a = 8'd29; b = 8'd86;  #10 
a = 8'd29; b = 8'd87;  #10 
a = 8'd29; b = 8'd88;  #10 
a = 8'd29; b = 8'd89;  #10 
a = 8'd29; b = 8'd90;  #10 
a = 8'd29; b = 8'd91;  #10 
a = 8'd29; b = 8'd92;  #10 
a = 8'd29; b = 8'd93;  #10 
a = 8'd29; b = 8'd94;  #10 
a = 8'd29; b = 8'd95;  #10 
a = 8'd29; b = 8'd96;  #10 
a = 8'd29; b = 8'd97;  #10 
a = 8'd29; b = 8'd98;  #10 
a = 8'd29; b = 8'd99;  #10 
a = 8'd29; b = 8'd100;  #10 
a = 8'd29; b = 8'd101;  #10 
a = 8'd29; b = 8'd102;  #10 
a = 8'd29; b = 8'd103;  #10 
a = 8'd29; b = 8'd104;  #10 
a = 8'd29; b = 8'd105;  #10 
a = 8'd29; b = 8'd106;  #10 
a = 8'd29; b = 8'd107;  #10 
a = 8'd29; b = 8'd108;  #10 
a = 8'd29; b = 8'd109;  #10 
a = 8'd29; b = 8'd110;  #10 
a = 8'd29; b = 8'd111;  #10 
a = 8'd29; b = 8'd112;  #10 
a = 8'd29; b = 8'd113;  #10 
a = 8'd29; b = 8'd114;  #10 
a = 8'd29; b = 8'd115;  #10 
a = 8'd29; b = 8'd116;  #10 
a = 8'd29; b = 8'd117;  #10 
a = 8'd29; b = 8'd118;  #10 
a = 8'd29; b = 8'd119;  #10 
a = 8'd29; b = 8'd120;  #10 
a = 8'd29; b = 8'd121;  #10 
a = 8'd29; b = 8'd122;  #10 
a = 8'd29; b = 8'd123;  #10 
a = 8'd29; b = 8'd124;  #10 
a = 8'd29; b = 8'd125;  #10 
a = 8'd29; b = 8'd126;  #10 
a = 8'd29; b = 8'd127;  #10 
a = 8'd29; b = 8'd128;  #10 
a = 8'd29; b = 8'd129;  #10 
a = 8'd29; b = 8'd130;  #10 
a = 8'd29; b = 8'd131;  #10 
a = 8'd29; b = 8'd132;  #10 
a = 8'd29; b = 8'd133;  #10 
a = 8'd29; b = 8'd134;  #10 
a = 8'd29; b = 8'd135;  #10 
a = 8'd29; b = 8'd136;  #10 
a = 8'd29; b = 8'd137;  #10 
a = 8'd29; b = 8'd138;  #10 
a = 8'd29; b = 8'd139;  #10 
a = 8'd29; b = 8'd140;  #10 
a = 8'd29; b = 8'd141;  #10 
a = 8'd29; b = 8'd142;  #10 
a = 8'd29; b = 8'd143;  #10 
a = 8'd29; b = 8'd144;  #10 
a = 8'd29; b = 8'd145;  #10 
a = 8'd29; b = 8'd146;  #10 
a = 8'd29; b = 8'd147;  #10 
a = 8'd29; b = 8'd148;  #10 
a = 8'd29; b = 8'd149;  #10 
a = 8'd29; b = 8'd150;  #10 
a = 8'd29; b = 8'd151;  #10 
a = 8'd29; b = 8'd152;  #10 
a = 8'd29; b = 8'd153;  #10 
a = 8'd29; b = 8'd154;  #10 
a = 8'd29; b = 8'd155;  #10 
a = 8'd29; b = 8'd156;  #10 
a = 8'd29; b = 8'd157;  #10 
a = 8'd29; b = 8'd158;  #10 
a = 8'd29; b = 8'd159;  #10 
a = 8'd29; b = 8'd160;  #10 
a = 8'd29; b = 8'd161;  #10 
a = 8'd29; b = 8'd162;  #10 
a = 8'd29; b = 8'd163;  #10 
a = 8'd29; b = 8'd164;  #10 
a = 8'd29; b = 8'd165;  #10 
a = 8'd29; b = 8'd166;  #10 
a = 8'd29; b = 8'd167;  #10 
a = 8'd29; b = 8'd168;  #10 
a = 8'd29; b = 8'd169;  #10 
a = 8'd29; b = 8'd170;  #10 
a = 8'd29; b = 8'd171;  #10 
a = 8'd29; b = 8'd172;  #10 
a = 8'd29; b = 8'd173;  #10 
a = 8'd29; b = 8'd174;  #10 
a = 8'd29; b = 8'd175;  #10 
a = 8'd29; b = 8'd176;  #10 
a = 8'd29; b = 8'd177;  #10 
a = 8'd29; b = 8'd178;  #10 
a = 8'd29; b = 8'd179;  #10 
a = 8'd29; b = 8'd180;  #10 
a = 8'd29; b = 8'd181;  #10 
a = 8'd29; b = 8'd182;  #10 
a = 8'd29; b = 8'd183;  #10 
a = 8'd29; b = 8'd184;  #10 
a = 8'd29; b = 8'd185;  #10 
a = 8'd29; b = 8'd186;  #10 
a = 8'd29; b = 8'd187;  #10 
a = 8'd29; b = 8'd188;  #10 
a = 8'd29; b = 8'd189;  #10 
a = 8'd29; b = 8'd190;  #10 
a = 8'd29; b = 8'd191;  #10 
a = 8'd29; b = 8'd192;  #10 
a = 8'd29; b = 8'd193;  #10 
a = 8'd29; b = 8'd194;  #10 
a = 8'd29; b = 8'd195;  #10 
a = 8'd29; b = 8'd196;  #10 
a = 8'd29; b = 8'd197;  #10 
a = 8'd29; b = 8'd198;  #10 
a = 8'd29; b = 8'd199;  #10 
a = 8'd29; b = 8'd200;  #10 
a = 8'd29; b = 8'd201;  #10 
a = 8'd29; b = 8'd202;  #10 
a = 8'd29; b = 8'd203;  #10 
a = 8'd29; b = 8'd204;  #10 
a = 8'd29; b = 8'd205;  #10 
a = 8'd29; b = 8'd206;  #10 
a = 8'd29; b = 8'd207;  #10 
a = 8'd29; b = 8'd208;  #10 
a = 8'd29; b = 8'd209;  #10 
a = 8'd29; b = 8'd210;  #10 
a = 8'd29; b = 8'd211;  #10 
a = 8'd29; b = 8'd212;  #10 
a = 8'd29; b = 8'd213;  #10 
a = 8'd29; b = 8'd214;  #10 
a = 8'd29; b = 8'd215;  #10 
a = 8'd29; b = 8'd216;  #10 
a = 8'd29; b = 8'd217;  #10 
a = 8'd29; b = 8'd218;  #10 
a = 8'd29; b = 8'd219;  #10 
a = 8'd29; b = 8'd220;  #10 
a = 8'd29; b = 8'd221;  #10 
a = 8'd29; b = 8'd222;  #10 
a = 8'd29; b = 8'd223;  #10 
a = 8'd29; b = 8'd224;  #10 
a = 8'd29; b = 8'd225;  #10 
a = 8'd29; b = 8'd226;  #10 
a = 8'd29; b = 8'd227;  #10 
a = 8'd29; b = 8'd228;  #10 
a = 8'd29; b = 8'd229;  #10 
a = 8'd29; b = 8'd230;  #10 
a = 8'd29; b = 8'd231;  #10 
a = 8'd29; b = 8'd232;  #10 
a = 8'd29; b = 8'd233;  #10 
a = 8'd29; b = 8'd234;  #10 
a = 8'd29; b = 8'd235;  #10 
a = 8'd29; b = 8'd236;  #10 
a = 8'd29; b = 8'd237;  #10 
a = 8'd29; b = 8'd238;  #10 
a = 8'd29; b = 8'd239;  #10 
a = 8'd29; b = 8'd240;  #10 
a = 8'd29; b = 8'd241;  #10 
a = 8'd29; b = 8'd242;  #10 
a = 8'd29; b = 8'd243;  #10 
a = 8'd29; b = 8'd244;  #10 
a = 8'd29; b = 8'd245;  #10 
a = 8'd29; b = 8'd246;  #10 
a = 8'd29; b = 8'd247;  #10 
a = 8'd29; b = 8'd248;  #10 
a = 8'd29; b = 8'd249;  #10 
a = 8'd29; b = 8'd250;  #10 
a = 8'd29; b = 8'd251;  #10 
a = 8'd29; b = 8'd252;  #10 
a = 8'd29; b = 8'd253;  #10 
a = 8'd29; b = 8'd254;  #10 
a = 8'd29; b = 8'd255;  #10 
a = 8'd30; b = 8'd0;  #10 
a = 8'd30; b = 8'd1;  #10 
a = 8'd30; b = 8'd2;  #10 
a = 8'd30; b = 8'd3;  #10 
a = 8'd30; b = 8'd4;  #10 
a = 8'd30; b = 8'd5;  #10 
a = 8'd30; b = 8'd6;  #10 
a = 8'd30; b = 8'd7;  #10 
a = 8'd30; b = 8'd8;  #10 
a = 8'd30; b = 8'd9;  #10 
a = 8'd30; b = 8'd10;  #10 
a = 8'd30; b = 8'd11;  #10 
a = 8'd30; b = 8'd12;  #10 
a = 8'd30; b = 8'd13;  #10 
a = 8'd30; b = 8'd14;  #10 
a = 8'd30; b = 8'd15;  #10 
a = 8'd30; b = 8'd16;  #10 
a = 8'd30; b = 8'd17;  #10 
a = 8'd30; b = 8'd18;  #10 
a = 8'd30; b = 8'd19;  #10 
a = 8'd30; b = 8'd20;  #10 
a = 8'd30; b = 8'd21;  #10 
a = 8'd30; b = 8'd22;  #10 
a = 8'd30; b = 8'd23;  #10 
a = 8'd30; b = 8'd24;  #10 
a = 8'd30; b = 8'd25;  #10 
a = 8'd30; b = 8'd26;  #10 
a = 8'd30; b = 8'd27;  #10 
a = 8'd30; b = 8'd28;  #10 
a = 8'd30; b = 8'd29;  #10 
a = 8'd30; b = 8'd30;  #10 
a = 8'd30; b = 8'd31;  #10 
a = 8'd30; b = 8'd32;  #10 
a = 8'd30; b = 8'd33;  #10 
a = 8'd30; b = 8'd34;  #10 
a = 8'd30; b = 8'd35;  #10 
a = 8'd30; b = 8'd36;  #10 
a = 8'd30; b = 8'd37;  #10 
a = 8'd30; b = 8'd38;  #10 
a = 8'd30; b = 8'd39;  #10 
a = 8'd30; b = 8'd40;  #10 
a = 8'd30; b = 8'd41;  #10 
a = 8'd30; b = 8'd42;  #10 
a = 8'd30; b = 8'd43;  #10 
a = 8'd30; b = 8'd44;  #10 
a = 8'd30; b = 8'd45;  #10 
a = 8'd30; b = 8'd46;  #10 
a = 8'd30; b = 8'd47;  #10 
a = 8'd30; b = 8'd48;  #10 
a = 8'd30; b = 8'd49;  #10 
a = 8'd30; b = 8'd50;  #10 
a = 8'd30; b = 8'd51;  #10 
a = 8'd30; b = 8'd52;  #10 
a = 8'd30; b = 8'd53;  #10 
a = 8'd30; b = 8'd54;  #10 
a = 8'd30; b = 8'd55;  #10 
a = 8'd30; b = 8'd56;  #10 
a = 8'd30; b = 8'd57;  #10 
a = 8'd30; b = 8'd58;  #10 
a = 8'd30; b = 8'd59;  #10 
a = 8'd30; b = 8'd60;  #10 
a = 8'd30; b = 8'd61;  #10 
a = 8'd30; b = 8'd62;  #10 
a = 8'd30; b = 8'd63;  #10 
a = 8'd30; b = 8'd64;  #10 
a = 8'd30; b = 8'd65;  #10 
a = 8'd30; b = 8'd66;  #10 
a = 8'd30; b = 8'd67;  #10 
a = 8'd30; b = 8'd68;  #10 
a = 8'd30; b = 8'd69;  #10 
a = 8'd30; b = 8'd70;  #10 
a = 8'd30; b = 8'd71;  #10 
a = 8'd30; b = 8'd72;  #10 
a = 8'd30; b = 8'd73;  #10 
a = 8'd30; b = 8'd74;  #10 
a = 8'd30; b = 8'd75;  #10 
a = 8'd30; b = 8'd76;  #10 
a = 8'd30; b = 8'd77;  #10 
a = 8'd30; b = 8'd78;  #10 
a = 8'd30; b = 8'd79;  #10 
a = 8'd30; b = 8'd80;  #10 
a = 8'd30; b = 8'd81;  #10 
a = 8'd30; b = 8'd82;  #10 
a = 8'd30; b = 8'd83;  #10 
a = 8'd30; b = 8'd84;  #10 
a = 8'd30; b = 8'd85;  #10 
a = 8'd30; b = 8'd86;  #10 
a = 8'd30; b = 8'd87;  #10 
a = 8'd30; b = 8'd88;  #10 
a = 8'd30; b = 8'd89;  #10 
a = 8'd30; b = 8'd90;  #10 
a = 8'd30; b = 8'd91;  #10 
a = 8'd30; b = 8'd92;  #10 
a = 8'd30; b = 8'd93;  #10 
a = 8'd30; b = 8'd94;  #10 
a = 8'd30; b = 8'd95;  #10 
a = 8'd30; b = 8'd96;  #10 
a = 8'd30; b = 8'd97;  #10 
a = 8'd30; b = 8'd98;  #10 
a = 8'd30; b = 8'd99;  #10 
a = 8'd30; b = 8'd100;  #10 
a = 8'd30; b = 8'd101;  #10 
a = 8'd30; b = 8'd102;  #10 
a = 8'd30; b = 8'd103;  #10 
a = 8'd30; b = 8'd104;  #10 
a = 8'd30; b = 8'd105;  #10 
a = 8'd30; b = 8'd106;  #10 
a = 8'd30; b = 8'd107;  #10 
a = 8'd30; b = 8'd108;  #10 
a = 8'd30; b = 8'd109;  #10 
a = 8'd30; b = 8'd110;  #10 
a = 8'd30; b = 8'd111;  #10 
a = 8'd30; b = 8'd112;  #10 
a = 8'd30; b = 8'd113;  #10 
a = 8'd30; b = 8'd114;  #10 
a = 8'd30; b = 8'd115;  #10 
a = 8'd30; b = 8'd116;  #10 
a = 8'd30; b = 8'd117;  #10 
a = 8'd30; b = 8'd118;  #10 
a = 8'd30; b = 8'd119;  #10 
a = 8'd30; b = 8'd120;  #10 
a = 8'd30; b = 8'd121;  #10 
a = 8'd30; b = 8'd122;  #10 
a = 8'd30; b = 8'd123;  #10 
a = 8'd30; b = 8'd124;  #10 
a = 8'd30; b = 8'd125;  #10 
a = 8'd30; b = 8'd126;  #10 
a = 8'd30; b = 8'd127;  #10 
a = 8'd30; b = 8'd128;  #10 
a = 8'd30; b = 8'd129;  #10 
a = 8'd30; b = 8'd130;  #10 
a = 8'd30; b = 8'd131;  #10 
a = 8'd30; b = 8'd132;  #10 
a = 8'd30; b = 8'd133;  #10 
a = 8'd30; b = 8'd134;  #10 
a = 8'd30; b = 8'd135;  #10 
a = 8'd30; b = 8'd136;  #10 
a = 8'd30; b = 8'd137;  #10 
a = 8'd30; b = 8'd138;  #10 
a = 8'd30; b = 8'd139;  #10 
a = 8'd30; b = 8'd140;  #10 
a = 8'd30; b = 8'd141;  #10 
a = 8'd30; b = 8'd142;  #10 
a = 8'd30; b = 8'd143;  #10 
a = 8'd30; b = 8'd144;  #10 
a = 8'd30; b = 8'd145;  #10 
a = 8'd30; b = 8'd146;  #10 
a = 8'd30; b = 8'd147;  #10 
a = 8'd30; b = 8'd148;  #10 
a = 8'd30; b = 8'd149;  #10 
a = 8'd30; b = 8'd150;  #10 
a = 8'd30; b = 8'd151;  #10 
a = 8'd30; b = 8'd152;  #10 
a = 8'd30; b = 8'd153;  #10 
a = 8'd30; b = 8'd154;  #10 
a = 8'd30; b = 8'd155;  #10 
a = 8'd30; b = 8'd156;  #10 
a = 8'd30; b = 8'd157;  #10 
a = 8'd30; b = 8'd158;  #10 
a = 8'd30; b = 8'd159;  #10 
a = 8'd30; b = 8'd160;  #10 
a = 8'd30; b = 8'd161;  #10 
a = 8'd30; b = 8'd162;  #10 
a = 8'd30; b = 8'd163;  #10 
a = 8'd30; b = 8'd164;  #10 
a = 8'd30; b = 8'd165;  #10 
a = 8'd30; b = 8'd166;  #10 
a = 8'd30; b = 8'd167;  #10 
a = 8'd30; b = 8'd168;  #10 
a = 8'd30; b = 8'd169;  #10 
a = 8'd30; b = 8'd170;  #10 
a = 8'd30; b = 8'd171;  #10 
a = 8'd30; b = 8'd172;  #10 
a = 8'd30; b = 8'd173;  #10 
a = 8'd30; b = 8'd174;  #10 
a = 8'd30; b = 8'd175;  #10 
a = 8'd30; b = 8'd176;  #10 
a = 8'd30; b = 8'd177;  #10 
a = 8'd30; b = 8'd178;  #10 
a = 8'd30; b = 8'd179;  #10 
a = 8'd30; b = 8'd180;  #10 
a = 8'd30; b = 8'd181;  #10 
a = 8'd30; b = 8'd182;  #10 
a = 8'd30; b = 8'd183;  #10 
a = 8'd30; b = 8'd184;  #10 
a = 8'd30; b = 8'd185;  #10 
a = 8'd30; b = 8'd186;  #10 
a = 8'd30; b = 8'd187;  #10 
a = 8'd30; b = 8'd188;  #10 
a = 8'd30; b = 8'd189;  #10 
a = 8'd30; b = 8'd190;  #10 
a = 8'd30; b = 8'd191;  #10 
a = 8'd30; b = 8'd192;  #10 
a = 8'd30; b = 8'd193;  #10 
a = 8'd30; b = 8'd194;  #10 
a = 8'd30; b = 8'd195;  #10 
a = 8'd30; b = 8'd196;  #10 
a = 8'd30; b = 8'd197;  #10 
a = 8'd30; b = 8'd198;  #10 
a = 8'd30; b = 8'd199;  #10 
a = 8'd30; b = 8'd200;  #10 
a = 8'd30; b = 8'd201;  #10 
a = 8'd30; b = 8'd202;  #10 
a = 8'd30; b = 8'd203;  #10 
a = 8'd30; b = 8'd204;  #10 
a = 8'd30; b = 8'd205;  #10 
a = 8'd30; b = 8'd206;  #10 
a = 8'd30; b = 8'd207;  #10 
a = 8'd30; b = 8'd208;  #10 
a = 8'd30; b = 8'd209;  #10 
a = 8'd30; b = 8'd210;  #10 
a = 8'd30; b = 8'd211;  #10 
a = 8'd30; b = 8'd212;  #10 
a = 8'd30; b = 8'd213;  #10 
a = 8'd30; b = 8'd214;  #10 
a = 8'd30; b = 8'd215;  #10 
a = 8'd30; b = 8'd216;  #10 
a = 8'd30; b = 8'd217;  #10 
a = 8'd30; b = 8'd218;  #10 
a = 8'd30; b = 8'd219;  #10 
a = 8'd30; b = 8'd220;  #10 
a = 8'd30; b = 8'd221;  #10 
a = 8'd30; b = 8'd222;  #10 
a = 8'd30; b = 8'd223;  #10 
a = 8'd30; b = 8'd224;  #10 
a = 8'd30; b = 8'd225;  #10 
a = 8'd30; b = 8'd226;  #10 
a = 8'd30; b = 8'd227;  #10 
a = 8'd30; b = 8'd228;  #10 
a = 8'd30; b = 8'd229;  #10 
a = 8'd30; b = 8'd230;  #10 
a = 8'd30; b = 8'd231;  #10 
a = 8'd30; b = 8'd232;  #10 
a = 8'd30; b = 8'd233;  #10 
a = 8'd30; b = 8'd234;  #10 
a = 8'd30; b = 8'd235;  #10 
a = 8'd30; b = 8'd236;  #10 
a = 8'd30; b = 8'd237;  #10 
a = 8'd30; b = 8'd238;  #10 
a = 8'd30; b = 8'd239;  #10 
a = 8'd30; b = 8'd240;  #10 
a = 8'd30; b = 8'd241;  #10 
a = 8'd30; b = 8'd242;  #10 
a = 8'd30; b = 8'd243;  #10 
a = 8'd30; b = 8'd244;  #10 
a = 8'd30; b = 8'd245;  #10 
a = 8'd30; b = 8'd246;  #10 
a = 8'd30; b = 8'd247;  #10 
a = 8'd30; b = 8'd248;  #10 
a = 8'd30; b = 8'd249;  #10 
a = 8'd30; b = 8'd250;  #10 
a = 8'd30; b = 8'd251;  #10 
a = 8'd30; b = 8'd252;  #10 
a = 8'd30; b = 8'd253;  #10 
a = 8'd30; b = 8'd254;  #10 
a = 8'd30; b = 8'd255;  #10 
a = 8'd31; b = 8'd0;  #10 
a = 8'd31; b = 8'd1;  #10 
a = 8'd31; b = 8'd2;  #10 
a = 8'd31; b = 8'd3;  #10 
a = 8'd31; b = 8'd4;  #10 
a = 8'd31; b = 8'd5;  #10 
a = 8'd31; b = 8'd6;  #10 
a = 8'd31; b = 8'd7;  #10 
a = 8'd31; b = 8'd8;  #10 
a = 8'd31; b = 8'd9;  #10 
a = 8'd31; b = 8'd10;  #10 
a = 8'd31; b = 8'd11;  #10 
a = 8'd31; b = 8'd12;  #10 
a = 8'd31; b = 8'd13;  #10 
a = 8'd31; b = 8'd14;  #10 
a = 8'd31; b = 8'd15;  #10 
a = 8'd31; b = 8'd16;  #10 
a = 8'd31; b = 8'd17;  #10 
a = 8'd31; b = 8'd18;  #10 
a = 8'd31; b = 8'd19;  #10 
a = 8'd31; b = 8'd20;  #10 
a = 8'd31; b = 8'd21;  #10 
a = 8'd31; b = 8'd22;  #10 
a = 8'd31; b = 8'd23;  #10 
a = 8'd31; b = 8'd24;  #10 
a = 8'd31; b = 8'd25;  #10 
a = 8'd31; b = 8'd26;  #10 
a = 8'd31; b = 8'd27;  #10 
a = 8'd31; b = 8'd28;  #10 
a = 8'd31; b = 8'd29;  #10 
a = 8'd31; b = 8'd30;  #10 
a = 8'd31; b = 8'd31;  #10 
a = 8'd31; b = 8'd32;  #10 
a = 8'd31; b = 8'd33;  #10 
a = 8'd31; b = 8'd34;  #10 
a = 8'd31; b = 8'd35;  #10 
a = 8'd31; b = 8'd36;  #10 
a = 8'd31; b = 8'd37;  #10 
a = 8'd31; b = 8'd38;  #10 
a = 8'd31; b = 8'd39;  #10 
a = 8'd31; b = 8'd40;  #10 
a = 8'd31; b = 8'd41;  #10 
a = 8'd31; b = 8'd42;  #10 
a = 8'd31; b = 8'd43;  #10 
a = 8'd31; b = 8'd44;  #10 
a = 8'd31; b = 8'd45;  #10 
a = 8'd31; b = 8'd46;  #10 
a = 8'd31; b = 8'd47;  #10 
a = 8'd31; b = 8'd48;  #10 
a = 8'd31; b = 8'd49;  #10 
a = 8'd31; b = 8'd50;  #10 
a = 8'd31; b = 8'd51;  #10 
a = 8'd31; b = 8'd52;  #10 
a = 8'd31; b = 8'd53;  #10 
a = 8'd31; b = 8'd54;  #10 
a = 8'd31; b = 8'd55;  #10 
a = 8'd31; b = 8'd56;  #10 
a = 8'd31; b = 8'd57;  #10 
a = 8'd31; b = 8'd58;  #10 
a = 8'd31; b = 8'd59;  #10 
a = 8'd31; b = 8'd60;  #10 
a = 8'd31; b = 8'd61;  #10 
a = 8'd31; b = 8'd62;  #10 
a = 8'd31; b = 8'd63;  #10 
a = 8'd31; b = 8'd64;  #10 
a = 8'd31; b = 8'd65;  #10 
a = 8'd31; b = 8'd66;  #10 
a = 8'd31; b = 8'd67;  #10 
a = 8'd31; b = 8'd68;  #10 
a = 8'd31; b = 8'd69;  #10 
a = 8'd31; b = 8'd70;  #10 
a = 8'd31; b = 8'd71;  #10 
a = 8'd31; b = 8'd72;  #10 
a = 8'd31; b = 8'd73;  #10 
a = 8'd31; b = 8'd74;  #10 
a = 8'd31; b = 8'd75;  #10 
a = 8'd31; b = 8'd76;  #10 
a = 8'd31; b = 8'd77;  #10 
a = 8'd31; b = 8'd78;  #10 
a = 8'd31; b = 8'd79;  #10 
a = 8'd31; b = 8'd80;  #10 
a = 8'd31; b = 8'd81;  #10 
a = 8'd31; b = 8'd82;  #10 
a = 8'd31; b = 8'd83;  #10 
a = 8'd31; b = 8'd84;  #10 
a = 8'd31; b = 8'd85;  #10 
a = 8'd31; b = 8'd86;  #10 
a = 8'd31; b = 8'd87;  #10 
a = 8'd31; b = 8'd88;  #10 
a = 8'd31; b = 8'd89;  #10 
a = 8'd31; b = 8'd90;  #10 
a = 8'd31; b = 8'd91;  #10 
a = 8'd31; b = 8'd92;  #10 
a = 8'd31; b = 8'd93;  #10 
a = 8'd31; b = 8'd94;  #10 
a = 8'd31; b = 8'd95;  #10 
a = 8'd31; b = 8'd96;  #10 
a = 8'd31; b = 8'd97;  #10 
a = 8'd31; b = 8'd98;  #10 
a = 8'd31; b = 8'd99;  #10 
a = 8'd31; b = 8'd100;  #10 
a = 8'd31; b = 8'd101;  #10 
a = 8'd31; b = 8'd102;  #10 
a = 8'd31; b = 8'd103;  #10 
a = 8'd31; b = 8'd104;  #10 
a = 8'd31; b = 8'd105;  #10 
a = 8'd31; b = 8'd106;  #10 
a = 8'd31; b = 8'd107;  #10 
a = 8'd31; b = 8'd108;  #10 
a = 8'd31; b = 8'd109;  #10 
a = 8'd31; b = 8'd110;  #10 
a = 8'd31; b = 8'd111;  #10 
a = 8'd31; b = 8'd112;  #10 
a = 8'd31; b = 8'd113;  #10 
a = 8'd31; b = 8'd114;  #10 
a = 8'd31; b = 8'd115;  #10 
a = 8'd31; b = 8'd116;  #10 
a = 8'd31; b = 8'd117;  #10 
a = 8'd31; b = 8'd118;  #10 
a = 8'd31; b = 8'd119;  #10 
a = 8'd31; b = 8'd120;  #10 
a = 8'd31; b = 8'd121;  #10 
a = 8'd31; b = 8'd122;  #10 
a = 8'd31; b = 8'd123;  #10 
a = 8'd31; b = 8'd124;  #10 
a = 8'd31; b = 8'd125;  #10 
a = 8'd31; b = 8'd126;  #10 
a = 8'd31; b = 8'd127;  #10 
a = 8'd31; b = 8'd128;  #10 
a = 8'd31; b = 8'd129;  #10 
a = 8'd31; b = 8'd130;  #10 
a = 8'd31; b = 8'd131;  #10 
a = 8'd31; b = 8'd132;  #10 
a = 8'd31; b = 8'd133;  #10 
a = 8'd31; b = 8'd134;  #10 
a = 8'd31; b = 8'd135;  #10 
a = 8'd31; b = 8'd136;  #10 
a = 8'd31; b = 8'd137;  #10 
a = 8'd31; b = 8'd138;  #10 
a = 8'd31; b = 8'd139;  #10 
a = 8'd31; b = 8'd140;  #10 
a = 8'd31; b = 8'd141;  #10 
a = 8'd31; b = 8'd142;  #10 
a = 8'd31; b = 8'd143;  #10 
a = 8'd31; b = 8'd144;  #10 
a = 8'd31; b = 8'd145;  #10 
a = 8'd31; b = 8'd146;  #10 
a = 8'd31; b = 8'd147;  #10 
a = 8'd31; b = 8'd148;  #10 
a = 8'd31; b = 8'd149;  #10 
a = 8'd31; b = 8'd150;  #10 
a = 8'd31; b = 8'd151;  #10 
a = 8'd31; b = 8'd152;  #10 
a = 8'd31; b = 8'd153;  #10 
a = 8'd31; b = 8'd154;  #10 
a = 8'd31; b = 8'd155;  #10 
a = 8'd31; b = 8'd156;  #10 
a = 8'd31; b = 8'd157;  #10 
a = 8'd31; b = 8'd158;  #10 
a = 8'd31; b = 8'd159;  #10 
a = 8'd31; b = 8'd160;  #10 
a = 8'd31; b = 8'd161;  #10 
a = 8'd31; b = 8'd162;  #10 
a = 8'd31; b = 8'd163;  #10 
a = 8'd31; b = 8'd164;  #10 
a = 8'd31; b = 8'd165;  #10 
a = 8'd31; b = 8'd166;  #10 
a = 8'd31; b = 8'd167;  #10 
a = 8'd31; b = 8'd168;  #10 
a = 8'd31; b = 8'd169;  #10 
a = 8'd31; b = 8'd170;  #10 
a = 8'd31; b = 8'd171;  #10 
a = 8'd31; b = 8'd172;  #10 
a = 8'd31; b = 8'd173;  #10 
a = 8'd31; b = 8'd174;  #10 
a = 8'd31; b = 8'd175;  #10 
a = 8'd31; b = 8'd176;  #10 
a = 8'd31; b = 8'd177;  #10 
a = 8'd31; b = 8'd178;  #10 
a = 8'd31; b = 8'd179;  #10 
a = 8'd31; b = 8'd180;  #10 
a = 8'd31; b = 8'd181;  #10 
a = 8'd31; b = 8'd182;  #10 
a = 8'd31; b = 8'd183;  #10 
a = 8'd31; b = 8'd184;  #10 
a = 8'd31; b = 8'd185;  #10 
a = 8'd31; b = 8'd186;  #10 
a = 8'd31; b = 8'd187;  #10 
a = 8'd31; b = 8'd188;  #10 
a = 8'd31; b = 8'd189;  #10 
a = 8'd31; b = 8'd190;  #10 
a = 8'd31; b = 8'd191;  #10 
a = 8'd31; b = 8'd192;  #10 
a = 8'd31; b = 8'd193;  #10 
a = 8'd31; b = 8'd194;  #10 
a = 8'd31; b = 8'd195;  #10 
a = 8'd31; b = 8'd196;  #10 
a = 8'd31; b = 8'd197;  #10 
a = 8'd31; b = 8'd198;  #10 
a = 8'd31; b = 8'd199;  #10 
a = 8'd31; b = 8'd200;  #10 
a = 8'd31; b = 8'd201;  #10 
a = 8'd31; b = 8'd202;  #10 
a = 8'd31; b = 8'd203;  #10 
a = 8'd31; b = 8'd204;  #10 
a = 8'd31; b = 8'd205;  #10 
a = 8'd31; b = 8'd206;  #10 
a = 8'd31; b = 8'd207;  #10 
a = 8'd31; b = 8'd208;  #10 
a = 8'd31; b = 8'd209;  #10 
a = 8'd31; b = 8'd210;  #10 
a = 8'd31; b = 8'd211;  #10 
a = 8'd31; b = 8'd212;  #10 
a = 8'd31; b = 8'd213;  #10 
a = 8'd31; b = 8'd214;  #10 
a = 8'd31; b = 8'd215;  #10 
a = 8'd31; b = 8'd216;  #10 
a = 8'd31; b = 8'd217;  #10 
a = 8'd31; b = 8'd218;  #10 
a = 8'd31; b = 8'd219;  #10 
a = 8'd31; b = 8'd220;  #10 
a = 8'd31; b = 8'd221;  #10 
a = 8'd31; b = 8'd222;  #10 
a = 8'd31; b = 8'd223;  #10 
a = 8'd31; b = 8'd224;  #10 
a = 8'd31; b = 8'd225;  #10 
a = 8'd31; b = 8'd226;  #10 
a = 8'd31; b = 8'd227;  #10 
a = 8'd31; b = 8'd228;  #10 
a = 8'd31; b = 8'd229;  #10 
a = 8'd31; b = 8'd230;  #10 
a = 8'd31; b = 8'd231;  #10 
a = 8'd31; b = 8'd232;  #10 
a = 8'd31; b = 8'd233;  #10 
a = 8'd31; b = 8'd234;  #10 
a = 8'd31; b = 8'd235;  #10 
a = 8'd31; b = 8'd236;  #10 
a = 8'd31; b = 8'd237;  #10 
a = 8'd31; b = 8'd238;  #10 
a = 8'd31; b = 8'd239;  #10 
a = 8'd31; b = 8'd240;  #10 
a = 8'd31; b = 8'd241;  #10 
a = 8'd31; b = 8'd242;  #10 
a = 8'd31; b = 8'd243;  #10 
a = 8'd31; b = 8'd244;  #10 
a = 8'd31; b = 8'd245;  #10 
a = 8'd31; b = 8'd246;  #10 
a = 8'd31; b = 8'd247;  #10 
a = 8'd31; b = 8'd248;  #10 
a = 8'd31; b = 8'd249;  #10 
a = 8'd31; b = 8'd250;  #10 
a = 8'd31; b = 8'd251;  #10 
a = 8'd31; b = 8'd252;  #10 
a = 8'd31; b = 8'd253;  #10 
a = 8'd31; b = 8'd254;  #10 
a = 8'd31; b = 8'd255;  #10 
a = 8'd32; b = 8'd0;  #10 
a = 8'd32; b = 8'd1;  #10 
a = 8'd32; b = 8'd2;  #10 
a = 8'd32; b = 8'd3;  #10 
a = 8'd32; b = 8'd4;  #10 
a = 8'd32; b = 8'd5;  #10 
a = 8'd32; b = 8'd6;  #10 
a = 8'd32; b = 8'd7;  #10 
a = 8'd32; b = 8'd8;  #10 
a = 8'd32; b = 8'd9;  #10 
a = 8'd32; b = 8'd10;  #10 
a = 8'd32; b = 8'd11;  #10 
a = 8'd32; b = 8'd12;  #10 
a = 8'd32; b = 8'd13;  #10 
a = 8'd32; b = 8'd14;  #10 
a = 8'd32; b = 8'd15;  #10 
a = 8'd32; b = 8'd16;  #10 
a = 8'd32; b = 8'd17;  #10 
a = 8'd32; b = 8'd18;  #10 
a = 8'd32; b = 8'd19;  #10 
a = 8'd32; b = 8'd20;  #10 
a = 8'd32; b = 8'd21;  #10 
a = 8'd32; b = 8'd22;  #10 
a = 8'd32; b = 8'd23;  #10 
a = 8'd32; b = 8'd24;  #10 
a = 8'd32; b = 8'd25;  #10 
a = 8'd32; b = 8'd26;  #10 
a = 8'd32; b = 8'd27;  #10 
a = 8'd32; b = 8'd28;  #10 
a = 8'd32; b = 8'd29;  #10 
a = 8'd32; b = 8'd30;  #10 
a = 8'd32; b = 8'd31;  #10 
a = 8'd32; b = 8'd32;  #10 
a = 8'd32; b = 8'd33;  #10 
a = 8'd32; b = 8'd34;  #10 
a = 8'd32; b = 8'd35;  #10 
a = 8'd32; b = 8'd36;  #10 
a = 8'd32; b = 8'd37;  #10 
a = 8'd32; b = 8'd38;  #10 
a = 8'd32; b = 8'd39;  #10 
a = 8'd32; b = 8'd40;  #10 
a = 8'd32; b = 8'd41;  #10 
a = 8'd32; b = 8'd42;  #10 
a = 8'd32; b = 8'd43;  #10 
a = 8'd32; b = 8'd44;  #10 
a = 8'd32; b = 8'd45;  #10 
a = 8'd32; b = 8'd46;  #10 
a = 8'd32; b = 8'd47;  #10 
a = 8'd32; b = 8'd48;  #10 
a = 8'd32; b = 8'd49;  #10 
a = 8'd32; b = 8'd50;  #10 
a = 8'd32; b = 8'd51;  #10 
a = 8'd32; b = 8'd52;  #10 
a = 8'd32; b = 8'd53;  #10 
a = 8'd32; b = 8'd54;  #10 
a = 8'd32; b = 8'd55;  #10 
a = 8'd32; b = 8'd56;  #10 
a = 8'd32; b = 8'd57;  #10 
a = 8'd32; b = 8'd58;  #10 
a = 8'd32; b = 8'd59;  #10 
a = 8'd32; b = 8'd60;  #10 
a = 8'd32; b = 8'd61;  #10 
a = 8'd32; b = 8'd62;  #10 
a = 8'd32; b = 8'd63;  #10 
a = 8'd32; b = 8'd64;  #10 
a = 8'd32; b = 8'd65;  #10 
a = 8'd32; b = 8'd66;  #10 
a = 8'd32; b = 8'd67;  #10 
a = 8'd32; b = 8'd68;  #10 
a = 8'd32; b = 8'd69;  #10 
a = 8'd32; b = 8'd70;  #10 
a = 8'd32; b = 8'd71;  #10 
a = 8'd32; b = 8'd72;  #10 
a = 8'd32; b = 8'd73;  #10 
a = 8'd32; b = 8'd74;  #10 
a = 8'd32; b = 8'd75;  #10 
a = 8'd32; b = 8'd76;  #10 
a = 8'd32; b = 8'd77;  #10 
a = 8'd32; b = 8'd78;  #10 
a = 8'd32; b = 8'd79;  #10 
a = 8'd32; b = 8'd80;  #10 
a = 8'd32; b = 8'd81;  #10 
a = 8'd32; b = 8'd82;  #10 
a = 8'd32; b = 8'd83;  #10 
a = 8'd32; b = 8'd84;  #10 
a = 8'd32; b = 8'd85;  #10 
a = 8'd32; b = 8'd86;  #10 
a = 8'd32; b = 8'd87;  #10 
a = 8'd32; b = 8'd88;  #10 
a = 8'd32; b = 8'd89;  #10 
a = 8'd32; b = 8'd90;  #10 
a = 8'd32; b = 8'd91;  #10 
a = 8'd32; b = 8'd92;  #10 
a = 8'd32; b = 8'd93;  #10 
a = 8'd32; b = 8'd94;  #10 
a = 8'd32; b = 8'd95;  #10 
a = 8'd32; b = 8'd96;  #10 
a = 8'd32; b = 8'd97;  #10 
a = 8'd32; b = 8'd98;  #10 
a = 8'd32; b = 8'd99;  #10 
a = 8'd32; b = 8'd100;  #10 
a = 8'd32; b = 8'd101;  #10 
a = 8'd32; b = 8'd102;  #10 
a = 8'd32; b = 8'd103;  #10 
a = 8'd32; b = 8'd104;  #10 
a = 8'd32; b = 8'd105;  #10 
a = 8'd32; b = 8'd106;  #10 
a = 8'd32; b = 8'd107;  #10 
a = 8'd32; b = 8'd108;  #10 
a = 8'd32; b = 8'd109;  #10 
a = 8'd32; b = 8'd110;  #10 
a = 8'd32; b = 8'd111;  #10 
a = 8'd32; b = 8'd112;  #10 
a = 8'd32; b = 8'd113;  #10 
a = 8'd32; b = 8'd114;  #10 
a = 8'd32; b = 8'd115;  #10 
a = 8'd32; b = 8'd116;  #10 
a = 8'd32; b = 8'd117;  #10 
a = 8'd32; b = 8'd118;  #10 
a = 8'd32; b = 8'd119;  #10 
a = 8'd32; b = 8'd120;  #10 
a = 8'd32; b = 8'd121;  #10 
a = 8'd32; b = 8'd122;  #10 
a = 8'd32; b = 8'd123;  #10 
a = 8'd32; b = 8'd124;  #10 
a = 8'd32; b = 8'd125;  #10 
a = 8'd32; b = 8'd126;  #10 
a = 8'd32; b = 8'd127;  #10 
a = 8'd32; b = 8'd128;  #10 
a = 8'd32; b = 8'd129;  #10 
a = 8'd32; b = 8'd130;  #10 
a = 8'd32; b = 8'd131;  #10 
a = 8'd32; b = 8'd132;  #10 
a = 8'd32; b = 8'd133;  #10 
a = 8'd32; b = 8'd134;  #10 
a = 8'd32; b = 8'd135;  #10 
a = 8'd32; b = 8'd136;  #10 
a = 8'd32; b = 8'd137;  #10 
a = 8'd32; b = 8'd138;  #10 
a = 8'd32; b = 8'd139;  #10 
a = 8'd32; b = 8'd140;  #10 
a = 8'd32; b = 8'd141;  #10 
a = 8'd32; b = 8'd142;  #10 
a = 8'd32; b = 8'd143;  #10 
a = 8'd32; b = 8'd144;  #10 
a = 8'd32; b = 8'd145;  #10 
a = 8'd32; b = 8'd146;  #10 
a = 8'd32; b = 8'd147;  #10 
a = 8'd32; b = 8'd148;  #10 
a = 8'd32; b = 8'd149;  #10 
a = 8'd32; b = 8'd150;  #10 
a = 8'd32; b = 8'd151;  #10 
a = 8'd32; b = 8'd152;  #10 
a = 8'd32; b = 8'd153;  #10 
a = 8'd32; b = 8'd154;  #10 
a = 8'd32; b = 8'd155;  #10 
a = 8'd32; b = 8'd156;  #10 
a = 8'd32; b = 8'd157;  #10 
a = 8'd32; b = 8'd158;  #10 
a = 8'd32; b = 8'd159;  #10 
a = 8'd32; b = 8'd160;  #10 
a = 8'd32; b = 8'd161;  #10 
a = 8'd32; b = 8'd162;  #10 
a = 8'd32; b = 8'd163;  #10 
a = 8'd32; b = 8'd164;  #10 
a = 8'd32; b = 8'd165;  #10 
a = 8'd32; b = 8'd166;  #10 
a = 8'd32; b = 8'd167;  #10 
a = 8'd32; b = 8'd168;  #10 
a = 8'd32; b = 8'd169;  #10 
a = 8'd32; b = 8'd170;  #10 
a = 8'd32; b = 8'd171;  #10 
a = 8'd32; b = 8'd172;  #10 
a = 8'd32; b = 8'd173;  #10 
a = 8'd32; b = 8'd174;  #10 
a = 8'd32; b = 8'd175;  #10 
a = 8'd32; b = 8'd176;  #10 
a = 8'd32; b = 8'd177;  #10 
a = 8'd32; b = 8'd178;  #10 
a = 8'd32; b = 8'd179;  #10 
a = 8'd32; b = 8'd180;  #10 
a = 8'd32; b = 8'd181;  #10 
a = 8'd32; b = 8'd182;  #10 
a = 8'd32; b = 8'd183;  #10 
a = 8'd32; b = 8'd184;  #10 
a = 8'd32; b = 8'd185;  #10 
a = 8'd32; b = 8'd186;  #10 
a = 8'd32; b = 8'd187;  #10 
a = 8'd32; b = 8'd188;  #10 
a = 8'd32; b = 8'd189;  #10 
a = 8'd32; b = 8'd190;  #10 
a = 8'd32; b = 8'd191;  #10 
a = 8'd32; b = 8'd192;  #10 
a = 8'd32; b = 8'd193;  #10 
a = 8'd32; b = 8'd194;  #10 
a = 8'd32; b = 8'd195;  #10 
a = 8'd32; b = 8'd196;  #10 
a = 8'd32; b = 8'd197;  #10 
a = 8'd32; b = 8'd198;  #10 
a = 8'd32; b = 8'd199;  #10 
a = 8'd32; b = 8'd200;  #10 
a = 8'd32; b = 8'd201;  #10 
a = 8'd32; b = 8'd202;  #10 
a = 8'd32; b = 8'd203;  #10 
a = 8'd32; b = 8'd204;  #10 
a = 8'd32; b = 8'd205;  #10 
a = 8'd32; b = 8'd206;  #10 
a = 8'd32; b = 8'd207;  #10 
a = 8'd32; b = 8'd208;  #10 
a = 8'd32; b = 8'd209;  #10 
a = 8'd32; b = 8'd210;  #10 
a = 8'd32; b = 8'd211;  #10 
a = 8'd32; b = 8'd212;  #10 
a = 8'd32; b = 8'd213;  #10 
a = 8'd32; b = 8'd214;  #10 
a = 8'd32; b = 8'd215;  #10 
a = 8'd32; b = 8'd216;  #10 
a = 8'd32; b = 8'd217;  #10 
a = 8'd32; b = 8'd218;  #10 
a = 8'd32; b = 8'd219;  #10 
a = 8'd32; b = 8'd220;  #10 
a = 8'd32; b = 8'd221;  #10 
a = 8'd32; b = 8'd222;  #10 
a = 8'd32; b = 8'd223;  #10 
a = 8'd32; b = 8'd224;  #10 
a = 8'd32; b = 8'd225;  #10 
a = 8'd32; b = 8'd226;  #10 
a = 8'd32; b = 8'd227;  #10 
a = 8'd32; b = 8'd228;  #10 
a = 8'd32; b = 8'd229;  #10 
a = 8'd32; b = 8'd230;  #10 
a = 8'd32; b = 8'd231;  #10 
a = 8'd32; b = 8'd232;  #10 
a = 8'd32; b = 8'd233;  #10 
a = 8'd32; b = 8'd234;  #10 
a = 8'd32; b = 8'd235;  #10 
a = 8'd32; b = 8'd236;  #10 
a = 8'd32; b = 8'd237;  #10 
a = 8'd32; b = 8'd238;  #10 
a = 8'd32; b = 8'd239;  #10 
a = 8'd32; b = 8'd240;  #10 
a = 8'd32; b = 8'd241;  #10 
a = 8'd32; b = 8'd242;  #10 
a = 8'd32; b = 8'd243;  #10 
a = 8'd32; b = 8'd244;  #10 
a = 8'd32; b = 8'd245;  #10 
a = 8'd32; b = 8'd246;  #10 
a = 8'd32; b = 8'd247;  #10 
a = 8'd32; b = 8'd248;  #10 
a = 8'd32; b = 8'd249;  #10 
a = 8'd32; b = 8'd250;  #10 
a = 8'd32; b = 8'd251;  #10 
a = 8'd32; b = 8'd252;  #10 
a = 8'd32; b = 8'd253;  #10 
a = 8'd32; b = 8'd254;  #10 
a = 8'd32; b = 8'd255;  #10 
a = 8'd33; b = 8'd0;  #10 
a = 8'd33; b = 8'd1;  #10 
a = 8'd33; b = 8'd2;  #10 
a = 8'd33; b = 8'd3;  #10 
a = 8'd33; b = 8'd4;  #10 
a = 8'd33; b = 8'd5;  #10 
a = 8'd33; b = 8'd6;  #10 
a = 8'd33; b = 8'd7;  #10 
a = 8'd33; b = 8'd8;  #10 
a = 8'd33; b = 8'd9;  #10 
a = 8'd33; b = 8'd10;  #10 
a = 8'd33; b = 8'd11;  #10 
a = 8'd33; b = 8'd12;  #10 
a = 8'd33; b = 8'd13;  #10 
a = 8'd33; b = 8'd14;  #10 
a = 8'd33; b = 8'd15;  #10 
a = 8'd33; b = 8'd16;  #10 
a = 8'd33; b = 8'd17;  #10 
a = 8'd33; b = 8'd18;  #10 
a = 8'd33; b = 8'd19;  #10 
a = 8'd33; b = 8'd20;  #10 
a = 8'd33; b = 8'd21;  #10 
a = 8'd33; b = 8'd22;  #10 
a = 8'd33; b = 8'd23;  #10 
a = 8'd33; b = 8'd24;  #10 
a = 8'd33; b = 8'd25;  #10 
a = 8'd33; b = 8'd26;  #10 
a = 8'd33; b = 8'd27;  #10 
a = 8'd33; b = 8'd28;  #10 
a = 8'd33; b = 8'd29;  #10 
a = 8'd33; b = 8'd30;  #10 
a = 8'd33; b = 8'd31;  #10 
a = 8'd33; b = 8'd32;  #10 
a = 8'd33; b = 8'd33;  #10 
a = 8'd33; b = 8'd34;  #10 
a = 8'd33; b = 8'd35;  #10 
a = 8'd33; b = 8'd36;  #10 
a = 8'd33; b = 8'd37;  #10 
a = 8'd33; b = 8'd38;  #10 
a = 8'd33; b = 8'd39;  #10 
a = 8'd33; b = 8'd40;  #10 
a = 8'd33; b = 8'd41;  #10 
a = 8'd33; b = 8'd42;  #10 
a = 8'd33; b = 8'd43;  #10 
a = 8'd33; b = 8'd44;  #10 
a = 8'd33; b = 8'd45;  #10 
a = 8'd33; b = 8'd46;  #10 
a = 8'd33; b = 8'd47;  #10 
a = 8'd33; b = 8'd48;  #10 
a = 8'd33; b = 8'd49;  #10 
a = 8'd33; b = 8'd50;  #10 
a = 8'd33; b = 8'd51;  #10 
a = 8'd33; b = 8'd52;  #10 
a = 8'd33; b = 8'd53;  #10 
a = 8'd33; b = 8'd54;  #10 
a = 8'd33; b = 8'd55;  #10 
a = 8'd33; b = 8'd56;  #10 
a = 8'd33; b = 8'd57;  #10 
a = 8'd33; b = 8'd58;  #10 
a = 8'd33; b = 8'd59;  #10 
a = 8'd33; b = 8'd60;  #10 
a = 8'd33; b = 8'd61;  #10 
a = 8'd33; b = 8'd62;  #10 
a = 8'd33; b = 8'd63;  #10 
a = 8'd33; b = 8'd64;  #10 
a = 8'd33; b = 8'd65;  #10 
a = 8'd33; b = 8'd66;  #10 
a = 8'd33; b = 8'd67;  #10 
a = 8'd33; b = 8'd68;  #10 
a = 8'd33; b = 8'd69;  #10 
a = 8'd33; b = 8'd70;  #10 
a = 8'd33; b = 8'd71;  #10 
a = 8'd33; b = 8'd72;  #10 
a = 8'd33; b = 8'd73;  #10 
a = 8'd33; b = 8'd74;  #10 
a = 8'd33; b = 8'd75;  #10 
a = 8'd33; b = 8'd76;  #10 
a = 8'd33; b = 8'd77;  #10 
a = 8'd33; b = 8'd78;  #10 
a = 8'd33; b = 8'd79;  #10 
a = 8'd33; b = 8'd80;  #10 
a = 8'd33; b = 8'd81;  #10 
a = 8'd33; b = 8'd82;  #10 
a = 8'd33; b = 8'd83;  #10 
a = 8'd33; b = 8'd84;  #10 
a = 8'd33; b = 8'd85;  #10 
a = 8'd33; b = 8'd86;  #10 
a = 8'd33; b = 8'd87;  #10 
a = 8'd33; b = 8'd88;  #10 
a = 8'd33; b = 8'd89;  #10 
a = 8'd33; b = 8'd90;  #10 
a = 8'd33; b = 8'd91;  #10 
a = 8'd33; b = 8'd92;  #10 
a = 8'd33; b = 8'd93;  #10 
a = 8'd33; b = 8'd94;  #10 
a = 8'd33; b = 8'd95;  #10 
a = 8'd33; b = 8'd96;  #10 
a = 8'd33; b = 8'd97;  #10 
a = 8'd33; b = 8'd98;  #10 
a = 8'd33; b = 8'd99;  #10 
a = 8'd33; b = 8'd100;  #10 
a = 8'd33; b = 8'd101;  #10 
a = 8'd33; b = 8'd102;  #10 
a = 8'd33; b = 8'd103;  #10 
a = 8'd33; b = 8'd104;  #10 
a = 8'd33; b = 8'd105;  #10 
a = 8'd33; b = 8'd106;  #10 
a = 8'd33; b = 8'd107;  #10 
a = 8'd33; b = 8'd108;  #10 
a = 8'd33; b = 8'd109;  #10 
a = 8'd33; b = 8'd110;  #10 
a = 8'd33; b = 8'd111;  #10 
a = 8'd33; b = 8'd112;  #10 
a = 8'd33; b = 8'd113;  #10 
a = 8'd33; b = 8'd114;  #10 
a = 8'd33; b = 8'd115;  #10 
a = 8'd33; b = 8'd116;  #10 
a = 8'd33; b = 8'd117;  #10 
a = 8'd33; b = 8'd118;  #10 
a = 8'd33; b = 8'd119;  #10 
a = 8'd33; b = 8'd120;  #10 
a = 8'd33; b = 8'd121;  #10 
a = 8'd33; b = 8'd122;  #10 
a = 8'd33; b = 8'd123;  #10 
a = 8'd33; b = 8'd124;  #10 
a = 8'd33; b = 8'd125;  #10 
a = 8'd33; b = 8'd126;  #10 
a = 8'd33; b = 8'd127;  #10 
a = 8'd33; b = 8'd128;  #10 
a = 8'd33; b = 8'd129;  #10 
a = 8'd33; b = 8'd130;  #10 
a = 8'd33; b = 8'd131;  #10 
a = 8'd33; b = 8'd132;  #10 
a = 8'd33; b = 8'd133;  #10 
a = 8'd33; b = 8'd134;  #10 
a = 8'd33; b = 8'd135;  #10 
a = 8'd33; b = 8'd136;  #10 
a = 8'd33; b = 8'd137;  #10 
a = 8'd33; b = 8'd138;  #10 
a = 8'd33; b = 8'd139;  #10 
a = 8'd33; b = 8'd140;  #10 
a = 8'd33; b = 8'd141;  #10 
a = 8'd33; b = 8'd142;  #10 
a = 8'd33; b = 8'd143;  #10 
a = 8'd33; b = 8'd144;  #10 
a = 8'd33; b = 8'd145;  #10 
a = 8'd33; b = 8'd146;  #10 
a = 8'd33; b = 8'd147;  #10 
a = 8'd33; b = 8'd148;  #10 
a = 8'd33; b = 8'd149;  #10 
a = 8'd33; b = 8'd150;  #10 
a = 8'd33; b = 8'd151;  #10 
a = 8'd33; b = 8'd152;  #10 
a = 8'd33; b = 8'd153;  #10 
a = 8'd33; b = 8'd154;  #10 
a = 8'd33; b = 8'd155;  #10 
a = 8'd33; b = 8'd156;  #10 
a = 8'd33; b = 8'd157;  #10 
a = 8'd33; b = 8'd158;  #10 
a = 8'd33; b = 8'd159;  #10 
a = 8'd33; b = 8'd160;  #10 
a = 8'd33; b = 8'd161;  #10 
a = 8'd33; b = 8'd162;  #10 
a = 8'd33; b = 8'd163;  #10 
a = 8'd33; b = 8'd164;  #10 
a = 8'd33; b = 8'd165;  #10 
a = 8'd33; b = 8'd166;  #10 
a = 8'd33; b = 8'd167;  #10 
a = 8'd33; b = 8'd168;  #10 
a = 8'd33; b = 8'd169;  #10 
a = 8'd33; b = 8'd170;  #10 
a = 8'd33; b = 8'd171;  #10 
a = 8'd33; b = 8'd172;  #10 
a = 8'd33; b = 8'd173;  #10 
a = 8'd33; b = 8'd174;  #10 
a = 8'd33; b = 8'd175;  #10 
a = 8'd33; b = 8'd176;  #10 
a = 8'd33; b = 8'd177;  #10 
a = 8'd33; b = 8'd178;  #10 
a = 8'd33; b = 8'd179;  #10 
a = 8'd33; b = 8'd180;  #10 
a = 8'd33; b = 8'd181;  #10 
a = 8'd33; b = 8'd182;  #10 
a = 8'd33; b = 8'd183;  #10 
a = 8'd33; b = 8'd184;  #10 
a = 8'd33; b = 8'd185;  #10 
a = 8'd33; b = 8'd186;  #10 
a = 8'd33; b = 8'd187;  #10 
a = 8'd33; b = 8'd188;  #10 
a = 8'd33; b = 8'd189;  #10 
a = 8'd33; b = 8'd190;  #10 
a = 8'd33; b = 8'd191;  #10 
a = 8'd33; b = 8'd192;  #10 
a = 8'd33; b = 8'd193;  #10 
a = 8'd33; b = 8'd194;  #10 
a = 8'd33; b = 8'd195;  #10 
a = 8'd33; b = 8'd196;  #10 
a = 8'd33; b = 8'd197;  #10 
a = 8'd33; b = 8'd198;  #10 
a = 8'd33; b = 8'd199;  #10 
a = 8'd33; b = 8'd200;  #10 
a = 8'd33; b = 8'd201;  #10 
a = 8'd33; b = 8'd202;  #10 
a = 8'd33; b = 8'd203;  #10 
a = 8'd33; b = 8'd204;  #10 
a = 8'd33; b = 8'd205;  #10 
a = 8'd33; b = 8'd206;  #10 
a = 8'd33; b = 8'd207;  #10 
a = 8'd33; b = 8'd208;  #10 
a = 8'd33; b = 8'd209;  #10 
a = 8'd33; b = 8'd210;  #10 
a = 8'd33; b = 8'd211;  #10 
a = 8'd33; b = 8'd212;  #10 
a = 8'd33; b = 8'd213;  #10 
a = 8'd33; b = 8'd214;  #10 
a = 8'd33; b = 8'd215;  #10 
a = 8'd33; b = 8'd216;  #10 
a = 8'd33; b = 8'd217;  #10 
a = 8'd33; b = 8'd218;  #10 
a = 8'd33; b = 8'd219;  #10 
a = 8'd33; b = 8'd220;  #10 
a = 8'd33; b = 8'd221;  #10 
a = 8'd33; b = 8'd222;  #10 
a = 8'd33; b = 8'd223;  #10 
a = 8'd33; b = 8'd224;  #10 
a = 8'd33; b = 8'd225;  #10 
a = 8'd33; b = 8'd226;  #10 
a = 8'd33; b = 8'd227;  #10 
a = 8'd33; b = 8'd228;  #10 
a = 8'd33; b = 8'd229;  #10 
a = 8'd33; b = 8'd230;  #10 
a = 8'd33; b = 8'd231;  #10 
a = 8'd33; b = 8'd232;  #10 
a = 8'd33; b = 8'd233;  #10 
a = 8'd33; b = 8'd234;  #10 
a = 8'd33; b = 8'd235;  #10 
a = 8'd33; b = 8'd236;  #10 
a = 8'd33; b = 8'd237;  #10 
a = 8'd33; b = 8'd238;  #10 
a = 8'd33; b = 8'd239;  #10 
a = 8'd33; b = 8'd240;  #10 
a = 8'd33; b = 8'd241;  #10 
a = 8'd33; b = 8'd242;  #10 
a = 8'd33; b = 8'd243;  #10 
a = 8'd33; b = 8'd244;  #10 
a = 8'd33; b = 8'd245;  #10 
a = 8'd33; b = 8'd246;  #10 
a = 8'd33; b = 8'd247;  #10 
a = 8'd33; b = 8'd248;  #10 
a = 8'd33; b = 8'd249;  #10 
a = 8'd33; b = 8'd250;  #10 
a = 8'd33; b = 8'd251;  #10 
a = 8'd33; b = 8'd252;  #10 
a = 8'd33; b = 8'd253;  #10 
a = 8'd33; b = 8'd254;  #10 
a = 8'd33; b = 8'd255;  #10 
a = 8'd34; b = 8'd0;  #10 
a = 8'd34; b = 8'd1;  #10 
a = 8'd34; b = 8'd2;  #10 
a = 8'd34; b = 8'd3;  #10 
a = 8'd34; b = 8'd4;  #10 
a = 8'd34; b = 8'd5;  #10 
a = 8'd34; b = 8'd6;  #10 
a = 8'd34; b = 8'd7;  #10 
a = 8'd34; b = 8'd8;  #10 
a = 8'd34; b = 8'd9;  #10 
a = 8'd34; b = 8'd10;  #10 
a = 8'd34; b = 8'd11;  #10 
a = 8'd34; b = 8'd12;  #10 
a = 8'd34; b = 8'd13;  #10 
a = 8'd34; b = 8'd14;  #10 
a = 8'd34; b = 8'd15;  #10 
a = 8'd34; b = 8'd16;  #10 
a = 8'd34; b = 8'd17;  #10 
a = 8'd34; b = 8'd18;  #10 
a = 8'd34; b = 8'd19;  #10 
a = 8'd34; b = 8'd20;  #10 
a = 8'd34; b = 8'd21;  #10 
a = 8'd34; b = 8'd22;  #10 
a = 8'd34; b = 8'd23;  #10 
a = 8'd34; b = 8'd24;  #10 
a = 8'd34; b = 8'd25;  #10 
a = 8'd34; b = 8'd26;  #10 
a = 8'd34; b = 8'd27;  #10 
a = 8'd34; b = 8'd28;  #10 
a = 8'd34; b = 8'd29;  #10 
a = 8'd34; b = 8'd30;  #10 
a = 8'd34; b = 8'd31;  #10 
a = 8'd34; b = 8'd32;  #10 
a = 8'd34; b = 8'd33;  #10 
a = 8'd34; b = 8'd34;  #10 
a = 8'd34; b = 8'd35;  #10 
a = 8'd34; b = 8'd36;  #10 
a = 8'd34; b = 8'd37;  #10 
a = 8'd34; b = 8'd38;  #10 
a = 8'd34; b = 8'd39;  #10 
a = 8'd34; b = 8'd40;  #10 
a = 8'd34; b = 8'd41;  #10 
a = 8'd34; b = 8'd42;  #10 
a = 8'd34; b = 8'd43;  #10 
a = 8'd34; b = 8'd44;  #10 
a = 8'd34; b = 8'd45;  #10 
a = 8'd34; b = 8'd46;  #10 
a = 8'd34; b = 8'd47;  #10 
a = 8'd34; b = 8'd48;  #10 
a = 8'd34; b = 8'd49;  #10 
a = 8'd34; b = 8'd50;  #10 
a = 8'd34; b = 8'd51;  #10 
a = 8'd34; b = 8'd52;  #10 
a = 8'd34; b = 8'd53;  #10 
a = 8'd34; b = 8'd54;  #10 
a = 8'd34; b = 8'd55;  #10 
a = 8'd34; b = 8'd56;  #10 
a = 8'd34; b = 8'd57;  #10 
a = 8'd34; b = 8'd58;  #10 
a = 8'd34; b = 8'd59;  #10 
a = 8'd34; b = 8'd60;  #10 
a = 8'd34; b = 8'd61;  #10 
a = 8'd34; b = 8'd62;  #10 
a = 8'd34; b = 8'd63;  #10 
a = 8'd34; b = 8'd64;  #10 
a = 8'd34; b = 8'd65;  #10 
a = 8'd34; b = 8'd66;  #10 
a = 8'd34; b = 8'd67;  #10 
a = 8'd34; b = 8'd68;  #10 
a = 8'd34; b = 8'd69;  #10 
a = 8'd34; b = 8'd70;  #10 
a = 8'd34; b = 8'd71;  #10 
a = 8'd34; b = 8'd72;  #10 
a = 8'd34; b = 8'd73;  #10 
a = 8'd34; b = 8'd74;  #10 
a = 8'd34; b = 8'd75;  #10 
a = 8'd34; b = 8'd76;  #10 
a = 8'd34; b = 8'd77;  #10 
a = 8'd34; b = 8'd78;  #10 
a = 8'd34; b = 8'd79;  #10 
a = 8'd34; b = 8'd80;  #10 
a = 8'd34; b = 8'd81;  #10 
a = 8'd34; b = 8'd82;  #10 
a = 8'd34; b = 8'd83;  #10 
a = 8'd34; b = 8'd84;  #10 
a = 8'd34; b = 8'd85;  #10 
a = 8'd34; b = 8'd86;  #10 
a = 8'd34; b = 8'd87;  #10 
a = 8'd34; b = 8'd88;  #10 
a = 8'd34; b = 8'd89;  #10 
a = 8'd34; b = 8'd90;  #10 
a = 8'd34; b = 8'd91;  #10 
a = 8'd34; b = 8'd92;  #10 
a = 8'd34; b = 8'd93;  #10 
a = 8'd34; b = 8'd94;  #10 
a = 8'd34; b = 8'd95;  #10 
a = 8'd34; b = 8'd96;  #10 
a = 8'd34; b = 8'd97;  #10 
a = 8'd34; b = 8'd98;  #10 
a = 8'd34; b = 8'd99;  #10 
a = 8'd34; b = 8'd100;  #10 
a = 8'd34; b = 8'd101;  #10 
a = 8'd34; b = 8'd102;  #10 
a = 8'd34; b = 8'd103;  #10 
a = 8'd34; b = 8'd104;  #10 
a = 8'd34; b = 8'd105;  #10 
a = 8'd34; b = 8'd106;  #10 
a = 8'd34; b = 8'd107;  #10 
a = 8'd34; b = 8'd108;  #10 
a = 8'd34; b = 8'd109;  #10 
a = 8'd34; b = 8'd110;  #10 
a = 8'd34; b = 8'd111;  #10 
a = 8'd34; b = 8'd112;  #10 
a = 8'd34; b = 8'd113;  #10 
a = 8'd34; b = 8'd114;  #10 
a = 8'd34; b = 8'd115;  #10 
a = 8'd34; b = 8'd116;  #10 
a = 8'd34; b = 8'd117;  #10 
a = 8'd34; b = 8'd118;  #10 
a = 8'd34; b = 8'd119;  #10 
a = 8'd34; b = 8'd120;  #10 
a = 8'd34; b = 8'd121;  #10 
a = 8'd34; b = 8'd122;  #10 
a = 8'd34; b = 8'd123;  #10 
a = 8'd34; b = 8'd124;  #10 
a = 8'd34; b = 8'd125;  #10 
a = 8'd34; b = 8'd126;  #10 
a = 8'd34; b = 8'd127;  #10 
a = 8'd34; b = 8'd128;  #10 
a = 8'd34; b = 8'd129;  #10 
a = 8'd34; b = 8'd130;  #10 
a = 8'd34; b = 8'd131;  #10 
a = 8'd34; b = 8'd132;  #10 
a = 8'd34; b = 8'd133;  #10 
a = 8'd34; b = 8'd134;  #10 
a = 8'd34; b = 8'd135;  #10 
a = 8'd34; b = 8'd136;  #10 
a = 8'd34; b = 8'd137;  #10 
a = 8'd34; b = 8'd138;  #10 
a = 8'd34; b = 8'd139;  #10 
a = 8'd34; b = 8'd140;  #10 
a = 8'd34; b = 8'd141;  #10 
a = 8'd34; b = 8'd142;  #10 
a = 8'd34; b = 8'd143;  #10 
a = 8'd34; b = 8'd144;  #10 
a = 8'd34; b = 8'd145;  #10 
a = 8'd34; b = 8'd146;  #10 
a = 8'd34; b = 8'd147;  #10 
a = 8'd34; b = 8'd148;  #10 
a = 8'd34; b = 8'd149;  #10 
a = 8'd34; b = 8'd150;  #10 
a = 8'd34; b = 8'd151;  #10 
a = 8'd34; b = 8'd152;  #10 
a = 8'd34; b = 8'd153;  #10 
a = 8'd34; b = 8'd154;  #10 
a = 8'd34; b = 8'd155;  #10 
a = 8'd34; b = 8'd156;  #10 
a = 8'd34; b = 8'd157;  #10 
a = 8'd34; b = 8'd158;  #10 
a = 8'd34; b = 8'd159;  #10 
a = 8'd34; b = 8'd160;  #10 
a = 8'd34; b = 8'd161;  #10 
a = 8'd34; b = 8'd162;  #10 
a = 8'd34; b = 8'd163;  #10 
a = 8'd34; b = 8'd164;  #10 
a = 8'd34; b = 8'd165;  #10 
a = 8'd34; b = 8'd166;  #10 
a = 8'd34; b = 8'd167;  #10 
a = 8'd34; b = 8'd168;  #10 
a = 8'd34; b = 8'd169;  #10 
a = 8'd34; b = 8'd170;  #10 
a = 8'd34; b = 8'd171;  #10 
a = 8'd34; b = 8'd172;  #10 
a = 8'd34; b = 8'd173;  #10 
a = 8'd34; b = 8'd174;  #10 
a = 8'd34; b = 8'd175;  #10 
a = 8'd34; b = 8'd176;  #10 
a = 8'd34; b = 8'd177;  #10 
a = 8'd34; b = 8'd178;  #10 
a = 8'd34; b = 8'd179;  #10 
a = 8'd34; b = 8'd180;  #10 
a = 8'd34; b = 8'd181;  #10 
a = 8'd34; b = 8'd182;  #10 
a = 8'd34; b = 8'd183;  #10 
a = 8'd34; b = 8'd184;  #10 
a = 8'd34; b = 8'd185;  #10 
a = 8'd34; b = 8'd186;  #10 
a = 8'd34; b = 8'd187;  #10 
a = 8'd34; b = 8'd188;  #10 
a = 8'd34; b = 8'd189;  #10 
a = 8'd34; b = 8'd190;  #10 
a = 8'd34; b = 8'd191;  #10 
a = 8'd34; b = 8'd192;  #10 
a = 8'd34; b = 8'd193;  #10 
a = 8'd34; b = 8'd194;  #10 
a = 8'd34; b = 8'd195;  #10 
a = 8'd34; b = 8'd196;  #10 
a = 8'd34; b = 8'd197;  #10 
a = 8'd34; b = 8'd198;  #10 
a = 8'd34; b = 8'd199;  #10 
a = 8'd34; b = 8'd200;  #10 
a = 8'd34; b = 8'd201;  #10 
a = 8'd34; b = 8'd202;  #10 
a = 8'd34; b = 8'd203;  #10 
a = 8'd34; b = 8'd204;  #10 
a = 8'd34; b = 8'd205;  #10 
a = 8'd34; b = 8'd206;  #10 
a = 8'd34; b = 8'd207;  #10 
a = 8'd34; b = 8'd208;  #10 
a = 8'd34; b = 8'd209;  #10 
a = 8'd34; b = 8'd210;  #10 
a = 8'd34; b = 8'd211;  #10 
a = 8'd34; b = 8'd212;  #10 
a = 8'd34; b = 8'd213;  #10 
a = 8'd34; b = 8'd214;  #10 
a = 8'd34; b = 8'd215;  #10 
a = 8'd34; b = 8'd216;  #10 
a = 8'd34; b = 8'd217;  #10 
a = 8'd34; b = 8'd218;  #10 
a = 8'd34; b = 8'd219;  #10 
a = 8'd34; b = 8'd220;  #10 
a = 8'd34; b = 8'd221;  #10 
a = 8'd34; b = 8'd222;  #10 
a = 8'd34; b = 8'd223;  #10 
a = 8'd34; b = 8'd224;  #10 
a = 8'd34; b = 8'd225;  #10 
a = 8'd34; b = 8'd226;  #10 
a = 8'd34; b = 8'd227;  #10 
a = 8'd34; b = 8'd228;  #10 
a = 8'd34; b = 8'd229;  #10 
a = 8'd34; b = 8'd230;  #10 
a = 8'd34; b = 8'd231;  #10 
a = 8'd34; b = 8'd232;  #10 
a = 8'd34; b = 8'd233;  #10 
a = 8'd34; b = 8'd234;  #10 
a = 8'd34; b = 8'd235;  #10 
a = 8'd34; b = 8'd236;  #10 
a = 8'd34; b = 8'd237;  #10 
a = 8'd34; b = 8'd238;  #10 
a = 8'd34; b = 8'd239;  #10 
a = 8'd34; b = 8'd240;  #10 
a = 8'd34; b = 8'd241;  #10 
a = 8'd34; b = 8'd242;  #10 
a = 8'd34; b = 8'd243;  #10 
a = 8'd34; b = 8'd244;  #10 
a = 8'd34; b = 8'd245;  #10 
a = 8'd34; b = 8'd246;  #10 
a = 8'd34; b = 8'd247;  #10 
a = 8'd34; b = 8'd248;  #10 
a = 8'd34; b = 8'd249;  #10 
a = 8'd34; b = 8'd250;  #10 
a = 8'd34; b = 8'd251;  #10 
a = 8'd34; b = 8'd252;  #10 
a = 8'd34; b = 8'd253;  #10 
a = 8'd34; b = 8'd254;  #10 
a = 8'd34; b = 8'd255;  #10 
a = 8'd35; b = 8'd0;  #10 
a = 8'd35; b = 8'd1;  #10 
a = 8'd35; b = 8'd2;  #10 
a = 8'd35; b = 8'd3;  #10 
a = 8'd35; b = 8'd4;  #10 
a = 8'd35; b = 8'd5;  #10 
a = 8'd35; b = 8'd6;  #10 
a = 8'd35; b = 8'd7;  #10 
a = 8'd35; b = 8'd8;  #10 
a = 8'd35; b = 8'd9;  #10 
a = 8'd35; b = 8'd10;  #10 
a = 8'd35; b = 8'd11;  #10 
a = 8'd35; b = 8'd12;  #10 
a = 8'd35; b = 8'd13;  #10 
a = 8'd35; b = 8'd14;  #10 
a = 8'd35; b = 8'd15;  #10 
a = 8'd35; b = 8'd16;  #10 
a = 8'd35; b = 8'd17;  #10 
a = 8'd35; b = 8'd18;  #10 
a = 8'd35; b = 8'd19;  #10 
a = 8'd35; b = 8'd20;  #10 
a = 8'd35; b = 8'd21;  #10 
a = 8'd35; b = 8'd22;  #10 
a = 8'd35; b = 8'd23;  #10 
a = 8'd35; b = 8'd24;  #10 
a = 8'd35; b = 8'd25;  #10 
a = 8'd35; b = 8'd26;  #10 
a = 8'd35; b = 8'd27;  #10 
a = 8'd35; b = 8'd28;  #10 
a = 8'd35; b = 8'd29;  #10 
a = 8'd35; b = 8'd30;  #10 
a = 8'd35; b = 8'd31;  #10 
a = 8'd35; b = 8'd32;  #10 
a = 8'd35; b = 8'd33;  #10 
a = 8'd35; b = 8'd34;  #10 
a = 8'd35; b = 8'd35;  #10 
a = 8'd35; b = 8'd36;  #10 
a = 8'd35; b = 8'd37;  #10 
a = 8'd35; b = 8'd38;  #10 
a = 8'd35; b = 8'd39;  #10 
a = 8'd35; b = 8'd40;  #10 
a = 8'd35; b = 8'd41;  #10 
a = 8'd35; b = 8'd42;  #10 
a = 8'd35; b = 8'd43;  #10 
a = 8'd35; b = 8'd44;  #10 
a = 8'd35; b = 8'd45;  #10 
a = 8'd35; b = 8'd46;  #10 
a = 8'd35; b = 8'd47;  #10 
a = 8'd35; b = 8'd48;  #10 
a = 8'd35; b = 8'd49;  #10 
a = 8'd35; b = 8'd50;  #10 
a = 8'd35; b = 8'd51;  #10 
a = 8'd35; b = 8'd52;  #10 
a = 8'd35; b = 8'd53;  #10 
a = 8'd35; b = 8'd54;  #10 
a = 8'd35; b = 8'd55;  #10 
a = 8'd35; b = 8'd56;  #10 
a = 8'd35; b = 8'd57;  #10 
a = 8'd35; b = 8'd58;  #10 
a = 8'd35; b = 8'd59;  #10 
a = 8'd35; b = 8'd60;  #10 
a = 8'd35; b = 8'd61;  #10 
a = 8'd35; b = 8'd62;  #10 
a = 8'd35; b = 8'd63;  #10 
a = 8'd35; b = 8'd64;  #10 
a = 8'd35; b = 8'd65;  #10 
a = 8'd35; b = 8'd66;  #10 
a = 8'd35; b = 8'd67;  #10 
a = 8'd35; b = 8'd68;  #10 
a = 8'd35; b = 8'd69;  #10 
a = 8'd35; b = 8'd70;  #10 
a = 8'd35; b = 8'd71;  #10 
a = 8'd35; b = 8'd72;  #10 
a = 8'd35; b = 8'd73;  #10 
a = 8'd35; b = 8'd74;  #10 
a = 8'd35; b = 8'd75;  #10 
a = 8'd35; b = 8'd76;  #10 
a = 8'd35; b = 8'd77;  #10 
a = 8'd35; b = 8'd78;  #10 
a = 8'd35; b = 8'd79;  #10 
a = 8'd35; b = 8'd80;  #10 
a = 8'd35; b = 8'd81;  #10 
a = 8'd35; b = 8'd82;  #10 
a = 8'd35; b = 8'd83;  #10 
a = 8'd35; b = 8'd84;  #10 
a = 8'd35; b = 8'd85;  #10 
a = 8'd35; b = 8'd86;  #10 
a = 8'd35; b = 8'd87;  #10 
a = 8'd35; b = 8'd88;  #10 
a = 8'd35; b = 8'd89;  #10 
a = 8'd35; b = 8'd90;  #10 
a = 8'd35; b = 8'd91;  #10 
a = 8'd35; b = 8'd92;  #10 
a = 8'd35; b = 8'd93;  #10 
a = 8'd35; b = 8'd94;  #10 
a = 8'd35; b = 8'd95;  #10 
a = 8'd35; b = 8'd96;  #10 
a = 8'd35; b = 8'd97;  #10 
a = 8'd35; b = 8'd98;  #10 
a = 8'd35; b = 8'd99;  #10 
a = 8'd35; b = 8'd100;  #10 
a = 8'd35; b = 8'd101;  #10 
a = 8'd35; b = 8'd102;  #10 
a = 8'd35; b = 8'd103;  #10 
a = 8'd35; b = 8'd104;  #10 
a = 8'd35; b = 8'd105;  #10 
a = 8'd35; b = 8'd106;  #10 
a = 8'd35; b = 8'd107;  #10 
a = 8'd35; b = 8'd108;  #10 
a = 8'd35; b = 8'd109;  #10 
a = 8'd35; b = 8'd110;  #10 
a = 8'd35; b = 8'd111;  #10 
a = 8'd35; b = 8'd112;  #10 
a = 8'd35; b = 8'd113;  #10 
a = 8'd35; b = 8'd114;  #10 
a = 8'd35; b = 8'd115;  #10 
a = 8'd35; b = 8'd116;  #10 
a = 8'd35; b = 8'd117;  #10 
a = 8'd35; b = 8'd118;  #10 
a = 8'd35; b = 8'd119;  #10 
a = 8'd35; b = 8'd120;  #10 
a = 8'd35; b = 8'd121;  #10 
a = 8'd35; b = 8'd122;  #10 
a = 8'd35; b = 8'd123;  #10 
a = 8'd35; b = 8'd124;  #10 
a = 8'd35; b = 8'd125;  #10 
a = 8'd35; b = 8'd126;  #10 
a = 8'd35; b = 8'd127;  #10 
a = 8'd35; b = 8'd128;  #10 
a = 8'd35; b = 8'd129;  #10 
a = 8'd35; b = 8'd130;  #10 
a = 8'd35; b = 8'd131;  #10 
a = 8'd35; b = 8'd132;  #10 
a = 8'd35; b = 8'd133;  #10 
a = 8'd35; b = 8'd134;  #10 
a = 8'd35; b = 8'd135;  #10 
a = 8'd35; b = 8'd136;  #10 
a = 8'd35; b = 8'd137;  #10 
a = 8'd35; b = 8'd138;  #10 
a = 8'd35; b = 8'd139;  #10 
a = 8'd35; b = 8'd140;  #10 
a = 8'd35; b = 8'd141;  #10 
a = 8'd35; b = 8'd142;  #10 
a = 8'd35; b = 8'd143;  #10 
a = 8'd35; b = 8'd144;  #10 
a = 8'd35; b = 8'd145;  #10 
a = 8'd35; b = 8'd146;  #10 
a = 8'd35; b = 8'd147;  #10 
a = 8'd35; b = 8'd148;  #10 
a = 8'd35; b = 8'd149;  #10 
a = 8'd35; b = 8'd150;  #10 
a = 8'd35; b = 8'd151;  #10 
a = 8'd35; b = 8'd152;  #10 
a = 8'd35; b = 8'd153;  #10 
a = 8'd35; b = 8'd154;  #10 
a = 8'd35; b = 8'd155;  #10 
a = 8'd35; b = 8'd156;  #10 
a = 8'd35; b = 8'd157;  #10 
a = 8'd35; b = 8'd158;  #10 
a = 8'd35; b = 8'd159;  #10 
a = 8'd35; b = 8'd160;  #10 
a = 8'd35; b = 8'd161;  #10 
a = 8'd35; b = 8'd162;  #10 
a = 8'd35; b = 8'd163;  #10 
a = 8'd35; b = 8'd164;  #10 
a = 8'd35; b = 8'd165;  #10 
a = 8'd35; b = 8'd166;  #10 
a = 8'd35; b = 8'd167;  #10 
a = 8'd35; b = 8'd168;  #10 
a = 8'd35; b = 8'd169;  #10 
a = 8'd35; b = 8'd170;  #10 
a = 8'd35; b = 8'd171;  #10 
a = 8'd35; b = 8'd172;  #10 
a = 8'd35; b = 8'd173;  #10 
a = 8'd35; b = 8'd174;  #10 
a = 8'd35; b = 8'd175;  #10 
a = 8'd35; b = 8'd176;  #10 
a = 8'd35; b = 8'd177;  #10 
a = 8'd35; b = 8'd178;  #10 
a = 8'd35; b = 8'd179;  #10 
a = 8'd35; b = 8'd180;  #10 
a = 8'd35; b = 8'd181;  #10 
a = 8'd35; b = 8'd182;  #10 
a = 8'd35; b = 8'd183;  #10 
a = 8'd35; b = 8'd184;  #10 
a = 8'd35; b = 8'd185;  #10 
a = 8'd35; b = 8'd186;  #10 
a = 8'd35; b = 8'd187;  #10 
a = 8'd35; b = 8'd188;  #10 
a = 8'd35; b = 8'd189;  #10 
a = 8'd35; b = 8'd190;  #10 
a = 8'd35; b = 8'd191;  #10 
a = 8'd35; b = 8'd192;  #10 
a = 8'd35; b = 8'd193;  #10 
a = 8'd35; b = 8'd194;  #10 
a = 8'd35; b = 8'd195;  #10 
a = 8'd35; b = 8'd196;  #10 
a = 8'd35; b = 8'd197;  #10 
a = 8'd35; b = 8'd198;  #10 
a = 8'd35; b = 8'd199;  #10 
a = 8'd35; b = 8'd200;  #10 
a = 8'd35; b = 8'd201;  #10 
a = 8'd35; b = 8'd202;  #10 
a = 8'd35; b = 8'd203;  #10 
a = 8'd35; b = 8'd204;  #10 
a = 8'd35; b = 8'd205;  #10 
a = 8'd35; b = 8'd206;  #10 
a = 8'd35; b = 8'd207;  #10 
a = 8'd35; b = 8'd208;  #10 
a = 8'd35; b = 8'd209;  #10 
a = 8'd35; b = 8'd210;  #10 
a = 8'd35; b = 8'd211;  #10 
a = 8'd35; b = 8'd212;  #10 
a = 8'd35; b = 8'd213;  #10 
a = 8'd35; b = 8'd214;  #10 
a = 8'd35; b = 8'd215;  #10 
a = 8'd35; b = 8'd216;  #10 
a = 8'd35; b = 8'd217;  #10 
a = 8'd35; b = 8'd218;  #10 
a = 8'd35; b = 8'd219;  #10 
a = 8'd35; b = 8'd220;  #10 
a = 8'd35; b = 8'd221;  #10 
a = 8'd35; b = 8'd222;  #10 
a = 8'd35; b = 8'd223;  #10 
a = 8'd35; b = 8'd224;  #10 
a = 8'd35; b = 8'd225;  #10 
a = 8'd35; b = 8'd226;  #10 
a = 8'd35; b = 8'd227;  #10 
a = 8'd35; b = 8'd228;  #10 
a = 8'd35; b = 8'd229;  #10 
a = 8'd35; b = 8'd230;  #10 
a = 8'd35; b = 8'd231;  #10 
a = 8'd35; b = 8'd232;  #10 
a = 8'd35; b = 8'd233;  #10 
a = 8'd35; b = 8'd234;  #10 
a = 8'd35; b = 8'd235;  #10 
a = 8'd35; b = 8'd236;  #10 
a = 8'd35; b = 8'd237;  #10 
a = 8'd35; b = 8'd238;  #10 
a = 8'd35; b = 8'd239;  #10 
a = 8'd35; b = 8'd240;  #10 
a = 8'd35; b = 8'd241;  #10 
a = 8'd35; b = 8'd242;  #10 
a = 8'd35; b = 8'd243;  #10 
a = 8'd35; b = 8'd244;  #10 
a = 8'd35; b = 8'd245;  #10 
a = 8'd35; b = 8'd246;  #10 
a = 8'd35; b = 8'd247;  #10 
a = 8'd35; b = 8'd248;  #10 
a = 8'd35; b = 8'd249;  #10 
a = 8'd35; b = 8'd250;  #10 
a = 8'd35; b = 8'd251;  #10 
a = 8'd35; b = 8'd252;  #10 
a = 8'd35; b = 8'd253;  #10 
a = 8'd35; b = 8'd254;  #10 
a = 8'd35; b = 8'd255;  #10 
a = 8'd36; b = 8'd0;  #10 
a = 8'd36; b = 8'd1;  #10 
a = 8'd36; b = 8'd2;  #10 
a = 8'd36; b = 8'd3;  #10 
a = 8'd36; b = 8'd4;  #10 
a = 8'd36; b = 8'd5;  #10 
a = 8'd36; b = 8'd6;  #10 
a = 8'd36; b = 8'd7;  #10 
a = 8'd36; b = 8'd8;  #10 
a = 8'd36; b = 8'd9;  #10 
a = 8'd36; b = 8'd10;  #10 
a = 8'd36; b = 8'd11;  #10 
a = 8'd36; b = 8'd12;  #10 
a = 8'd36; b = 8'd13;  #10 
a = 8'd36; b = 8'd14;  #10 
a = 8'd36; b = 8'd15;  #10 
a = 8'd36; b = 8'd16;  #10 
a = 8'd36; b = 8'd17;  #10 
a = 8'd36; b = 8'd18;  #10 
a = 8'd36; b = 8'd19;  #10 
a = 8'd36; b = 8'd20;  #10 
a = 8'd36; b = 8'd21;  #10 
a = 8'd36; b = 8'd22;  #10 
a = 8'd36; b = 8'd23;  #10 
a = 8'd36; b = 8'd24;  #10 
a = 8'd36; b = 8'd25;  #10 
a = 8'd36; b = 8'd26;  #10 
a = 8'd36; b = 8'd27;  #10 
a = 8'd36; b = 8'd28;  #10 
a = 8'd36; b = 8'd29;  #10 
a = 8'd36; b = 8'd30;  #10 
a = 8'd36; b = 8'd31;  #10 
a = 8'd36; b = 8'd32;  #10 
a = 8'd36; b = 8'd33;  #10 
a = 8'd36; b = 8'd34;  #10 
a = 8'd36; b = 8'd35;  #10 
a = 8'd36; b = 8'd36;  #10 
a = 8'd36; b = 8'd37;  #10 
a = 8'd36; b = 8'd38;  #10 
a = 8'd36; b = 8'd39;  #10 
a = 8'd36; b = 8'd40;  #10 
a = 8'd36; b = 8'd41;  #10 
a = 8'd36; b = 8'd42;  #10 
a = 8'd36; b = 8'd43;  #10 
a = 8'd36; b = 8'd44;  #10 
a = 8'd36; b = 8'd45;  #10 
a = 8'd36; b = 8'd46;  #10 
a = 8'd36; b = 8'd47;  #10 
a = 8'd36; b = 8'd48;  #10 
a = 8'd36; b = 8'd49;  #10 
a = 8'd36; b = 8'd50;  #10 
a = 8'd36; b = 8'd51;  #10 
a = 8'd36; b = 8'd52;  #10 
a = 8'd36; b = 8'd53;  #10 
a = 8'd36; b = 8'd54;  #10 
a = 8'd36; b = 8'd55;  #10 
a = 8'd36; b = 8'd56;  #10 
a = 8'd36; b = 8'd57;  #10 
a = 8'd36; b = 8'd58;  #10 
a = 8'd36; b = 8'd59;  #10 
a = 8'd36; b = 8'd60;  #10 
a = 8'd36; b = 8'd61;  #10 
a = 8'd36; b = 8'd62;  #10 
a = 8'd36; b = 8'd63;  #10 
a = 8'd36; b = 8'd64;  #10 
a = 8'd36; b = 8'd65;  #10 
a = 8'd36; b = 8'd66;  #10 
a = 8'd36; b = 8'd67;  #10 
a = 8'd36; b = 8'd68;  #10 
a = 8'd36; b = 8'd69;  #10 
a = 8'd36; b = 8'd70;  #10 
a = 8'd36; b = 8'd71;  #10 
a = 8'd36; b = 8'd72;  #10 
a = 8'd36; b = 8'd73;  #10 
a = 8'd36; b = 8'd74;  #10 
a = 8'd36; b = 8'd75;  #10 
a = 8'd36; b = 8'd76;  #10 
a = 8'd36; b = 8'd77;  #10 
a = 8'd36; b = 8'd78;  #10 
a = 8'd36; b = 8'd79;  #10 
a = 8'd36; b = 8'd80;  #10 
a = 8'd36; b = 8'd81;  #10 
a = 8'd36; b = 8'd82;  #10 
a = 8'd36; b = 8'd83;  #10 
a = 8'd36; b = 8'd84;  #10 
a = 8'd36; b = 8'd85;  #10 
a = 8'd36; b = 8'd86;  #10 
a = 8'd36; b = 8'd87;  #10 
a = 8'd36; b = 8'd88;  #10 
a = 8'd36; b = 8'd89;  #10 
a = 8'd36; b = 8'd90;  #10 
a = 8'd36; b = 8'd91;  #10 
a = 8'd36; b = 8'd92;  #10 
a = 8'd36; b = 8'd93;  #10 
a = 8'd36; b = 8'd94;  #10 
a = 8'd36; b = 8'd95;  #10 
a = 8'd36; b = 8'd96;  #10 
a = 8'd36; b = 8'd97;  #10 
a = 8'd36; b = 8'd98;  #10 
a = 8'd36; b = 8'd99;  #10 
a = 8'd36; b = 8'd100;  #10 
a = 8'd36; b = 8'd101;  #10 
a = 8'd36; b = 8'd102;  #10 
a = 8'd36; b = 8'd103;  #10 
a = 8'd36; b = 8'd104;  #10 
a = 8'd36; b = 8'd105;  #10 
a = 8'd36; b = 8'd106;  #10 
a = 8'd36; b = 8'd107;  #10 
a = 8'd36; b = 8'd108;  #10 
a = 8'd36; b = 8'd109;  #10 
a = 8'd36; b = 8'd110;  #10 
a = 8'd36; b = 8'd111;  #10 
a = 8'd36; b = 8'd112;  #10 
a = 8'd36; b = 8'd113;  #10 
a = 8'd36; b = 8'd114;  #10 
a = 8'd36; b = 8'd115;  #10 
a = 8'd36; b = 8'd116;  #10 
a = 8'd36; b = 8'd117;  #10 
a = 8'd36; b = 8'd118;  #10 
a = 8'd36; b = 8'd119;  #10 
a = 8'd36; b = 8'd120;  #10 
a = 8'd36; b = 8'd121;  #10 
a = 8'd36; b = 8'd122;  #10 
a = 8'd36; b = 8'd123;  #10 
a = 8'd36; b = 8'd124;  #10 
a = 8'd36; b = 8'd125;  #10 
a = 8'd36; b = 8'd126;  #10 
a = 8'd36; b = 8'd127;  #10 
a = 8'd36; b = 8'd128;  #10 
a = 8'd36; b = 8'd129;  #10 
a = 8'd36; b = 8'd130;  #10 
a = 8'd36; b = 8'd131;  #10 
a = 8'd36; b = 8'd132;  #10 
a = 8'd36; b = 8'd133;  #10 
a = 8'd36; b = 8'd134;  #10 
a = 8'd36; b = 8'd135;  #10 
a = 8'd36; b = 8'd136;  #10 
a = 8'd36; b = 8'd137;  #10 
a = 8'd36; b = 8'd138;  #10 
a = 8'd36; b = 8'd139;  #10 
a = 8'd36; b = 8'd140;  #10 
a = 8'd36; b = 8'd141;  #10 
a = 8'd36; b = 8'd142;  #10 
a = 8'd36; b = 8'd143;  #10 
a = 8'd36; b = 8'd144;  #10 
a = 8'd36; b = 8'd145;  #10 
a = 8'd36; b = 8'd146;  #10 
a = 8'd36; b = 8'd147;  #10 
a = 8'd36; b = 8'd148;  #10 
a = 8'd36; b = 8'd149;  #10 
a = 8'd36; b = 8'd150;  #10 
a = 8'd36; b = 8'd151;  #10 
a = 8'd36; b = 8'd152;  #10 
a = 8'd36; b = 8'd153;  #10 
a = 8'd36; b = 8'd154;  #10 
a = 8'd36; b = 8'd155;  #10 
a = 8'd36; b = 8'd156;  #10 
a = 8'd36; b = 8'd157;  #10 
a = 8'd36; b = 8'd158;  #10 
a = 8'd36; b = 8'd159;  #10 
a = 8'd36; b = 8'd160;  #10 
a = 8'd36; b = 8'd161;  #10 
a = 8'd36; b = 8'd162;  #10 
a = 8'd36; b = 8'd163;  #10 
a = 8'd36; b = 8'd164;  #10 
a = 8'd36; b = 8'd165;  #10 
a = 8'd36; b = 8'd166;  #10 
a = 8'd36; b = 8'd167;  #10 
a = 8'd36; b = 8'd168;  #10 
a = 8'd36; b = 8'd169;  #10 
a = 8'd36; b = 8'd170;  #10 
a = 8'd36; b = 8'd171;  #10 
a = 8'd36; b = 8'd172;  #10 
a = 8'd36; b = 8'd173;  #10 
a = 8'd36; b = 8'd174;  #10 
a = 8'd36; b = 8'd175;  #10 
a = 8'd36; b = 8'd176;  #10 
a = 8'd36; b = 8'd177;  #10 
a = 8'd36; b = 8'd178;  #10 
a = 8'd36; b = 8'd179;  #10 
a = 8'd36; b = 8'd180;  #10 
a = 8'd36; b = 8'd181;  #10 
a = 8'd36; b = 8'd182;  #10 
a = 8'd36; b = 8'd183;  #10 
a = 8'd36; b = 8'd184;  #10 
a = 8'd36; b = 8'd185;  #10 
a = 8'd36; b = 8'd186;  #10 
a = 8'd36; b = 8'd187;  #10 
a = 8'd36; b = 8'd188;  #10 
a = 8'd36; b = 8'd189;  #10 
a = 8'd36; b = 8'd190;  #10 
a = 8'd36; b = 8'd191;  #10 
a = 8'd36; b = 8'd192;  #10 
a = 8'd36; b = 8'd193;  #10 
a = 8'd36; b = 8'd194;  #10 
a = 8'd36; b = 8'd195;  #10 
a = 8'd36; b = 8'd196;  #10 
a = 8'd36; b = 8'd197;  #10 
a = 8'd36; b = 8'd198;  #10 
a = 8'd36; b = 8'd199;  #10 
a = 8'd36; b = 8'd200;  #10 
a = 8'd36; b = 8'd201;  #10 
a = 8'd36; b = 8'd202;  #10 
a = 8'd36; b = 8'd203;  #10 
a = 8'd36; b = 8'd204;  #10 
a = 8'd36; b = 8'd205;  #10 
a = 8'd36; b = 8'd206;  #10 
a = 8'd36; b = 8'd207;  #10 
a = 8'd36; b = 8'd208;  #10 
a = 8'd36; b = 8'd209;  #10 
a = 8'd36; b = 8'd210;  #10 
a = 8'd36; b = 8'd211;  #10 
a = 8'd36; b = 8'd212;  #10 
a = 8'd36; b = 8'd213;  #10 
a = 8'd36; b = 8'd214;  #10 
a = 8'd36; b = 8'd215;  #10 
a = 8'd36; b = 8'd216;  #10 
a = 8'd36; b = 8'd217;  #10 
a = 8'd36; b = 8'd218;  #10 
a = 8'd36; b = 8'd219;  #10 
a = 8'd36; b = 8'd220;  #10 
a = 8'd36; b = 8'd221;  #10 
a = 8'd36; b = 8'd222;  #10 
a = 8'd36; b = 8'd223;  #10 
a = 8'd36; b = 8'd224;  #10 
a = 8'd36; b = 8'd225;  #10 
a = 8'd36; b = 8'd226;  #10 
a = 8'd36; b = 8'd227;  #10 
a = 8'd36; b = 8'd228;  #10 
a = 8'd36; b = 8'd229;  #10 
a = 8'd36; b = 8'd230;  #10 
a = 8'd36; b = 8'd231;  #10 
a = 8'd36; b = 8'd232;  #10 
a = 8'd36; b = 8'd233;  #10 
a = 8'd36; b = 8'd234;  #10 
a = 8'd36; b = 8'd235;  #10 
a = 8'd36; b = 8'd236;  #10 
a = 8'd36; b = 8'd237;  #10 
a = 8'd36; b = 8'd238;  #10 
a = 8'd36; b = 8'd239;  #10 
a = 8'd36; b = 8'd240;  #10 
a = 8'd36; b = 8'd241;  #10 
a = 8'd36; b = 8'd242;  #10 
a = 8'd36; b = 8'd243;  #10 
a = 8'd36; b = 8'd244;  #10 
a = 8'd36; b = 8'd245;  #10 
a = 8'd36; b = 8'd246;  #10 
a = 8'd36; b = 8'd247;  #10 
a = 8'd36; b = 8'd248;  #10 
a = 8'd36; b = 8'd249;  #10 
a = 8'd36; b = 8'd250;  #10 
a = 8'd36; b = 8'd251;  #10 
a = 8'd36; b = 8'd252;  #10 
a = 8'd36; b = 8'd253;  #10 
a = 8'd36; b = 8'd254;  #10 
a = 8'd36; b = 8'd255;  #10 
a = 8'd37; b = 8'd0;  #10 
a = 8'd37; b = 8'd1;  #10 
a = 8'd37; b = 8'd2;  #10 
a = 8'd37; b = 8'd3;  #10 
a = 8'd37; b = 8'd4;  #10 
a = 8'd37; b = 8'd5;  #10 
a = 8'd37; b = 8'd6;  #10 
a = 8'd37; b = 8'd7;  #10 
a = 8'd37; b = 8'd8;  #10 
a = 8'd37; b = 8'd9;  #10 
a = 8'd37; b = 8'd10;  #10 
a = 8'd37; b = 8'd11;  #10 
a = 8'd37; b = 8'd12;  #10 
a = 8'd37; b = 8'd13;  #10 
a = 8'd37; b = 8'd14;  #10 
a = 8'd37; b = 8'd15;  #10 
a = 8'd37; b = 8'd16;  #10 
a = 8'd37; b = 8'd17;  #10 
a = 8'd37; b = 8'd18;  #10 
a = 8'd37; b = 8'd19;  #10 
a = 8'd37; b = 8'd20;  #10 
a = 8'd37; b = 8'd21;  #10 
a = 8'd37; b = 8'd22;  #10 
a = 8'd37; b = 8'd23;  #10 
a = 8'd37; b = 8'd24;  #10 
a = 8'd37; b = 8'd25;  #10 
a = 8'd37; b = 8'd26;  #10 
a = 8'd37; b = 8'd27;  #10 
a = 8'd37; b = 8'd28;  #10 
a = 8'd37; b = 8'd29;  #10 
a = 8'd37; b = 8'd30;  #10 
a = 8'd37; b = 8'd31;  #10 
a = 8'd37; b = 8'd32;  #10 
a = 8'd37; b = 8'd33;  #10 
a = 8'd37; b = 8'd34;  #10 
a = 8'd37; b = 8'd35;  #10 
a = 8'd37; b = 8'd36;  #10 
a = 8'd37; b = 8'd37;  #10 
a = 8'd37; b = 8'd38;  #10 
a = 8'd37; b = 8'd39;  #10 
a = 8'd37; b = 8'd40;  #10 
a = 8'd37; b = 8'd41;  #10 
a = 8'd37; b = 8'd42;  #10 
a = 8'd37; b = 8'd43;  #10 
a = 8'd37; b = 8'd44;  #10 
a = 8'd37; b = 8'd45;  #10 
a = 8'd37; b = 8'd46;  #10 
a = 8'd37; b = 8'd47;  #10 
a = 8'd37; b = 8'd48;  #10 
a = 8'd37; b = 8'd49;  #10 
a = 8'd37; b = 8'd50;  #10 
a = 8'd37; b = 8'd51;  #10 
a = 8'd37; b = 8'd52;  #10 
a = 8'd37; b = 8'd53;  #10 
a = 8'd37; b = 8'd54;  #10 
a = 8'd37; b = 8'd55;  #10 
a = 8'd37; b = 8'd56;  #10 
a = 8'd37; b = 8'd57;  #10 
a = 8'd37; b = 8'd58;  #10 
a = 8'd37; b = 8'd59;  #10 
a = 8'd37; b = 8'd60;  #10 
a = 8'd37; b = 8'd61;  #10 
a = 8'd37; b = 8'd62;  #10 
a = 8'd37; b = 8'd63;  #10 
a = 8'd37; b = 8'd64;  #10 
a = 8'd37; b = 8'd65;  #10 
a = 8'd37; b = 8'd66;  #10 
a = 8'd37; b = 8'd67;  #10 
a = 8'd37; b = 8'd68;  #10 
a = 8'd37; b = 8'd69;  #10 
a = 8'd37; b = 8'd70;  #10 
a = 8'd37; b = 8'd71;  #10 
a = 8'd37; b = 8'd72;  #10 
a = 8'd37; b = 8'd73;  #10 
a = 8'd37; b = 8'd74;  #10 
a = 8'd37; b = 8'd75;  #10 
a = 8'd37; b = 8'd76;  #10 
a = 8'd37; b = 8'd77;  #10 
a = 8'd37; b = 8'd78;  #10 
a = 8'd37; b = 8'd79;  #10 
a = 8'd37; b = 8'd80;  #10 
a = 8'd37; b = 8'd81;  #10 
a = 8'd37; b = 8'd82;  #10 
a = 8'd37; b = 8'd83;  #10 
a = 8'd37; b = 8'd84;  #10 
a = 8'd37; b = 8'd85;  #10 
a = 8'd37; b = 8'd86;  #10 
a = 8'd37; b = 8'd87;  #10 
a = 8'd37; b = 8'd88;  #10 
a = 8'd37; b = 8'd89;  #10 
a = 8'd37; b = 8'd90;  #10 
a = 8'd37; b = 8'd91;  #10 
a = 8'd37; b = 8'd92;  #10 
a = 8'd37; b = 8'd93;  #10 
a = 8'd37; b = 8'd94;  #10 
a = 8'd37; b = 8'd95;  #10 
a = 8'd37; b = 8'd96;  #10 
a = 8'd37; b = 8'd97;  #10 
a = 8'd37; b = 8'd98;  #10 
a = 8'd37; b = 8'd99;  #10 
a = 8'd37; b = 8'd100;  #10 
a = 8'd37; b = 8'd101;  #10 
a = 8'd37; b = 8'd102;  #10 
a = 8'd37; b = 8'd103;  #10 
a = 8'd37; b = 8'd104;  #10 
a = 8'd37; b = 8'd105;  #10 
a = 8'd37; b = 8'd106;  #10 
a = 8'd37; b = 8'd107;  #10 
a = 8'd37; b = 8'd108;  #10 
a = 8'd37; b = 8'd109;  #10 
a = 8'd37; b = 8'd110;  #10 
a = 8'd37; b = 8'd111;  #10 
a = 8'd37; b = 8'd112;  #10 
a = 8'd37; b = 8'd113;  #10 
a = 8'd37; b = 8'd114;  #10 
a = 8'd37; b = 8'd115;  #10 
a = 8'd37; b = 8'd116;  #10 
a = 8'd37; b = 8'd117;  #10 
a = 8'd37; b = 8'd118;  #10 
a = 8'd37; b = 8'd119;  #10 
a = 8'd37; b = 8'd120;  #10 
a = 8'd37; b = 8'd121;  #10 
a = 8'd37; b = 8'd122;  #10 
a = 8'd37; b = 8'd123;  #10 
a = 8'd37; b = 8'd124;  #10 
a = 8'd37; b = 8'd125;  #10 
a = 8'd37; b = 8'd126;  #10 
a = 8'd37; b = 8'd127;  #10 
a = 8'd37; b = 8'd128;  #10 
a = 8'd37; b = 8'd129;  #10 
a = 8'd37; b = 8'd130;  #10 
a = 8'd37; b = 8'd131;  #10 
a = 8'd37; b = 8'd132;  #10 
a = 8'd37; b = 8'd133;  #10 
a = 8'd37; b = 8'd134;  #10 
a = 8'd37; b = 8'd135;  #10 
a = 8'd37; b = 8'd136;  #10 
a = 8'd37; b = 8'd137;  #10 
a = 8'd37; b = 8'd138;  #10 
a = 8'd37; b = 8'd139;  #10 
a = 8'd37; b = 8'd140;  #10 
a = 8'd37; b = 8'd141;  #10 
a = 8'd37; b = 8'd142;  #10 
a = 8'd37; b = 8'd143;  #10 
a = 8'd37; b = 8'd144;  #10 
a = 8'd37; b = 8'd145;  #10 
a = 8'd37; b = 8'd146;  #10 
a = 8'd37; b = 8'd147;  #10 
a = 8'd37; b = 8'd148;  #10 
a = 8'd37; b = 8'd149;  #10 
a = 8'd37; b = 8'd150;  #10 
a = 8'd37; b = 8'd151;  #10 
a = 8'd37; b = 8'd152;  #10 
a = 8'd37; b = 8'd153;  #10 
a = 8'd37; b = 8'd154;  #10 
a = 8'd37; b = 8'd155;  #10 
a = 8'd37; b = 8'd156;  #10 
a = 8'd37; b = 8'd157;  #10 
a = 8'd37; b = 8'd158;  #10 
a = 8'd37; b = 8'd159;  #10 
a = 8'd37; b = 8'd160;  #10 
a = 8'd37; b = 8'd161;  #10 
a = 8'd37; b = 8'd162;  #10 
a = 8'd37; b = 8'd163;  #10 
a = 8'd37; b = 8'd164;  #10 
a = 8'd37; b = 8'd165;  #10 
a = 8'd37; b = 8'd166;  #10 
a = 8'd37; b = 8'd167;  #10 
a = 8'd37; b = 8'd168;  #10 
a = 8'd37; b = 8'd169;  #10 
a = 8'd37; b = 8'd170;  #10 
a = 8'd37; b = 8'd171;  #10 
a = 8'd37; b = 8'd172;  #10 
a = 8'd37; b = 8'd173;  #10 
a = 8'd37; b = 8'd174;  #10 
a = 8'd37; b = 8'd175;  #10 
a = 8'd37; b = 8'd176;  #10 
a = 8'd37; b = 8'd177;  #10 
a = 8'd37; b = 8'd178;  #10 
a = 8'd37; b = 8'd179;  #10 
a = 8'd37; b = 8'd180;  #10 
a = 8'd37; b = 8'd181;  #10 
a = 8'd37; b = 8'd182;  #10 
a = 8'd37; b = 8'd183;  #10 
a = 8'd37; b = 8'd184;  #10 
a = 8'd37; b = 8'd185;  #10 
a = 8'd37; b = 8'd186;  #10 
a = 8'd37; b = 8'd187;  #10 
a = 8'd37; b = 8'd188;  #10 
a = 8'd37; b = 8'd189;  #10 
a = 8'd37; b = 8'd190;  #10 
a = 8'd37; b = 8'd191;  #10 
a = 8'd37; b = 8'd192;  #10 
a = 8'd37; b = 8'd193;  #10 
a = 8'd37; b = 8'd194;  #10 
a = 8'd37; b = 8'd195;  #10 
a = 8'd37; b = 8'd196;  #10 
a = 8'd37; b = 8'd197;  #10 
a = 8'd37; b = 8'd198;  #10 
a = 8'd37; b = 8'd199;  #10 
a = 8'd37; b = 8'd200;  #10 
a = 8'd37; b = 8'd201;  #10 
a = 8'd37; b = 8'd202;  #10 
a = 8'd37; b = 8'd203;  #10 
a = 8'd37; b = 8'd204;  #10 
a = 8'd37; b = 8'd205;  #10 
a = 8'd37; b = 8'd206;  #10 
a = 8'd37; b = 8'd207;  #10 
a = 8'd37; b = 8'd208;  #10 
a = 8'd37; b = 8'd209;  #10 
a = 8'd37; b = 8'd210;  #10 
a = 8'd37; b = 8'd211;  #10 
a = 8'd37; b = 8'd212;  #10 
a = 8'd37; b = 8'd213;  #10 
a = 8'd37; b = 8'd214;  #10 
a = 8'd37; b = 8'd215;  #10 
a = 8'd37; b = 8'd216;  #10 
a = 8'd37; b = 8'd217;  #10 
a = 8'd37; b = 8'd218;  #10 
a = 8'd37; b = 8'd219;  #10 
a = 8'd37; b = 8'd220;  #10 
a = 8'd37; b = 8'd221;  #10 
a = 8'd37; b = 8'd222;  #10 
a = 8'd37; b = 8'd223;  #10 
a = 8'd37; b = 8'd224;  #10 
a = 8'd37; b = 8'd225;  #10 
a = 8'd37; b = 8'd226;  #10 
a = 8'd37; b = 8'd227;  #10 
a = 8'd37; b = 8'd228;  #10 
a = 8'd37; b = 8'd229;  #10 
a = 8'd37; b = 8'd230;  #10 
a = 8'd37; b = 8'd231;  #10 
a = 8'd37; b = 8'd232;  #10 
a = 8'd37; b = 8'd233;  #10 
a = 8'd37; b = 8'd234;  #10 
a = 8'd37; b = 8'd235;  #10 
a = 8'd37; b = 8'd236;  #10 
a = 8'd37; b = 8'd237;  #10 
a = 8'd37; b = 8'd238;  #10 
a = 8'd37; b = 8'd239;  #10 
a = 8'd37; b = 8'd240;  #10 
a = 8'd37; b = 8'd241;  #10 
a = 8'd37; b = 8'd242;  #10 
a = 8'd37; b = 8'd243;  #10 
a = 8'd37; b = 8'd244;  #10 
a = 8'd37; b = 8'd245;  #10 
a = 8'd37; b = 8'd246;  #10 
a = 8'd37; b = 8'd247;  #10 
a = 8'd37; b = 8'd248;  #10 
a = 8'd37; b = 8'd249;  #10 
a = 8'd37; b = 8'd250;  #10 
a = 8'd37; b = 8'd251;  #10 
a = 8'd37; b = 8'd252;  #10 
a = 8'd37; b = 8'd253;  #10 
a = 8'd37; b = 8'd254;  #10 
a = 8'd37; b = 8'd255;  #10 
a = 8'd38; b = 8'd0;  #10 
a = 8'd38; b = 8'd1;  #10 
a = 8'd38; b = 8'd2;  #10 
a = 8'd38; b = 8'd3;  #10 
a = 8'd38; b = 8'd4;  #10 
a = 8'd38; b = 8'd5;  #10 
a = 8'd38; b = 8'd6;  #10 
a = 8'd38; b = 8'd7;  #10 
a = 8'd38; b = 8'd8;  #10 
a = 8'd38; b = 8'd9;  #10 
a = 8'd38; b = 8'd10;  #10 
a = 8'd38; b = 8'd11;  #10 
a = 8'd38; b = 8'd12;  #10 
a = 8'd38; b = 8'd13;  #10 
a = 8'd38; b = 8'd14;  #10 
a = 8'd38; b = 8'd15;  #10 
a = 8'd38; b = 8'd16;  #10 
a = 8'd38; b = 8'd17;  #10 
a = 8'd38; b = 8'd18;  #10 
a = 8'd38; b = 8'd19;  #10 
a = 8'd38; b = 8'd20;  #10 
a = 8'd38; b = 8'd21;  #10 
a = 8'd38; b = 8'd22;  #10 
a = 8'd38; b = 8'd23;  #10 
a = 8'd38; b = 8'd24;  #10 
a = 8'd38; b = 8'd25;  #10 
a = 8'd38; b = 8'd26;  #10 
a = 8'd38; b = 8'd27;  #10 
a = 8'd38; b = 8'd28;  #10 
a = 8'd38; b = 8'd29;  #10 
a = 8'd38; b = 8'd30;  #10 
a = 8'd38; b = 8'd31;  #10 
a = 8'd38; b = 8'd32;  #10 
a = 8'd38; b = 8'd33;  #10 
a = 8'd38; b = 8'd34;  #10 
a = 8'd38; b = 8'd35;  #10 
a = 8'd38; b = 8'd36;  #10 
a = 8'd38; b = 8'd37;  #10 
a = 8'd38; b = 8'd38;  #10 
a = 8'd38; b = 8'd39;  #10 
a = 8'd38; b = 8'd40;  #10 
a = 8'd38; b = 8'd41;  #10 
a = 8'd38; b = 8'd42;  #10 
a = 8'd38; b = 8'd43;  #10 
a = 8'd38; b = 8'd44;  #10 
a = 8'd38; b = 8'd45;  #10 
a = 8'd38; b = 8'd46;  #10 
a = 8'd38; b = 8'd47;  #10 
a = 8'd38; b = 8'd48;  #10 
a = 8'd38; b = 8'd49;  #10 
a = 8'd38; b = 8'd50;  #10 
a = 8'd38; b = 8'd51;  #10 
a = 8'd38; b = 8'd52;  #10 
a = 8'd38; b = 8'd53;  #10 
a = 8'd38; b = 8'd54;  #10 
a = 8'd38; b = 8'd55;  #10 
a = 8'd38; b = 8'd56;  #10 
a = 8'd38; b = 8'd57;  #10 
a = 8'd38; b = 8'd58;  #10 
a = 8'd38; b = 8'd59;  #10 
a = 8'd38; b = 8'd60;  #10 
a = 8'd38; b = 8'd61;  #10 
a = 8'd38; b = 8'd62;  #10 
a = 8'd38; b = 8'd63;  #10 
a = 8'd38; b = 8'd64;  #10 
a = 8'd38; b = 8'd65;  #10 
a = 8'd38; b = 8'd66;  #10 
a = 8'd38; b = 8'd67;  #10 
a = 8'd38; b = 8'd68;  #10 
a = 8'd38; b = 8'd69;  #10 
a = 8'd38; b = 8'd70;  #10 
a = 8'd38; b = 8'd71;  #10 
a = 8'd38; b = 8'd72;  #10 
a = 8'd38; b = 8'd73;  #10 
a = 8'd38; b = 8'd74;  #10 
a = 8'd38; b = 8'd75;  #10 
a = 8'd38; b = 8'd76;  #10 
a = 8'd38; b = 8'd77;  #10 
a = 8'd38; b = 8'd78;  #10 
a = 8'd38; b = 8'd79;  #10 
a = 8'd38; b = 8'd80;  #10 
a = 8'd38; b = 8'd81;  #10 
a = 8'd38; b = 8'd82;  #10 
a = 8'd38; b = 8'd83;  #10 
a = 8'd38; b = 8'd84;  #10 
a = 8'd38; b = 8'd85;  #10 
a = 8'd38; b = 8'd86;  #10 
a = 8'd38; b = 8'd87;  #10 
a = 8'd38; b = 8'd88;  #10 
a = 8'd38; b = 8'd89;  #10 
a = 8'd38; b = 8'd90;  #10 
a = 8'd38; b = 8'd91;  #10 
a = 8'd38; b = 8'd92;  #10 
a = 8'd38; b = 8'd93;  #10 
a = 8'd38; b = 8'd94;  #10 
a = 8'd38; b = 8'd95;  #10 
a = 8'd38; b = 8'd96;  #10 
a = 8'd38; b = 8'd97;  #10 
a = 8'd38; b = 8'd98;  #10 
a = 8'd38; b = 8'd99;  #10 
a = 8'd38; b = 8'd100;  #10 
a = 8'd38; b = 8'd101;  #10 
a = 8'd38; b = 8'd102;  #10 
a = 8'd38; b = 8'd103;  #10 
a = 8'd38; b = 8'd104;  #10 
a = 8'd38; b = 8'd105;  #10 
a = 8'd38; b = 8'd106;  #10 
a = 8'd38; b = 8'd107;  #10 
a = 8'd38; b = 8'd108;  #10 
a = 8'd38; b = 8'd109;  #10 
a = 8'd38; b = 8'd110;  #10 
a = 8'd38; b = 8'd111;  #10 
a = 8'd38; b = 8'd112;  #10 
a = 8'd38; b = 8'd113;  #10 
a = 8'd38; b = 8'd114;  #10 
a = 8'd38; b = 8'd115;  #10 
a = 8'd38; b = 8'd116;  #10 
a = 8'd38; b = 8'd117;  #10 
a = 8'd38; b = 8'd118;  #10 
a = 8'd38; b = 8'd119;  #10 
a = 8'd38; b = 8'd120;  #10 
a = 8'd38; b = 8'd121;  #10 
a = 8'd38; b = 8'd122;  #10 
a = 8'd38; b = 8'd123;  #10 
a = 8'd38; b = 8'd124;  #10 
a = 8'd38; b = 8'd125;  #10 
a = 8'd38; b = 8'd126;  #10 
a = 8'd38; b = 8'd127;  #10 
a = 8'd38; b = 8'd128;  #10 
a = 8'd38; b = 8'd129;  #10 
a = 8'd38; b = 8'd130;  #10 
a = 8'd38; b = 8'd131;  #10 
a = 8'd38; b = 8'd132;  #10 
a = 8'd38; b = 8'd133;  #10 
a = 8'd38; b = 8'd134;  #10 
a = 8'd38; b = 8'd135;  #10 
a = 8'd38; b = 8'd136;  #10 
a = 8'd38; b = 8'd137;  #10 
a = 8'd38; b = 8'd138;  #10 
a = 8'd38; b = 8'd139;  #10 
a = 8'd38; b = 8'd140;  #10 
a = 8'd38; b = 8'd141;  #10 
a = 8'd38; b = 8'd142;  #10 
a = 8'd38; b = 8'd143;  #10 
a = 8'd38; b = 8'd144;  #10 
a = 8'd38; b = 8'd145;  #10 
a = 8'd38; b = 8'd146;  #10 
a = 8'd38; b = 8'd147;  #10 
a = 8'd38; b = 8'd148;  #10 
a = 8'd38; b = 8'd149;  #10 
a = 8'd38; b = 8'd150;  #10 
a = 8'd38; b = 8'd151;  #10 
a = 8'd38; b = 8'd152;  #10 
a = 8'd38; b = 8'd153;  #10 
a = 8'd38; b = 8'd154;  #10 
a = 8'd38; b = 8'd155;  #10 
a = 8'd38; b = 8'd156;  #10 
a = 8'd38; b = 8'd157;  #10 
a = 8'd38; b = 8'd158;  #10 
a = 8'd38; b = 8'd159;  #10 
a = 8'd38; b = 8'd160;  #10 
a = 8'd38; b = 8'd161;  #10 
a = 8'd38; b = 8'd162;  #10 
a = 8'd38; b = 8'd163;  #10 
a = 8'd38; b = 8'd164;  #10 
a = 8'd38; b = 8'd165;  #10 
a = 8'd38; b = 8'd166;  #10 
a = 8'd38; b = 8'd167;  #10 
a = 8'd38; b = 8'd168;  #10 
a = 8'd38; b = 8'd169;  #10 
a = 8'd38; b = 8'd170;  #10 
a = 8'd38; b = 8'd171;  #10 
a = 8'd38; b = 8'd172;  #10 
a = 8'd38; b = 8'd173;  #10 
a = 8'd38; b = 8'd174;  #10 
a = 8'd38; b = 8'd175;  #10 
a = 8'd38; b = 8'd176;  #10 
a = 8'd38; b = 8'd177;  #10 
a = 8'd38; b = 8'd178;  #10 
a = 8'd38; b = 8'd179;  #10 
a = 8'd38; b = 8'd180;  #10 
a = 8'd38; b = 8'd181;  #10 
a = 8'd38; b = 8'd182;  #10 
a = 8'd38; b = 8'd183;  #10 
a = 8'd38; b = 8'd184;  #10 
a = 8'd38; b = 8'd185;  #10 
a = 8'd38; b = 8'd186;  #10 
a = 8'd38; b = 8'd187;  #10 
a = 8'd38; b = 8'd188;  #10 
a = 8'd38; b = 8'd189;  #10 
a = 8'd38; b = 8'd190;  #10 
a = 8'd38; b = 8'd191;  #10 
a = 8'd38; b = 8'd192;  #10 
a = 8'd38; b = 8'd193;  #10 
a = 8'd38; b = 8'd194;  #10 
a = 8'd38; b = 8'd195;  #10 
a = 8'd38; b = 8'd196;  #10 
a = 8'd38; b = 8'd197;  #10 
a = 8'd38; b = 8'd198;  #10 
a = 8'd38; b = 8'd199;  #10 
a = 8'd38; b = 8'd200;  #10 
a = 8'd38; b = 8'd201;  #10 
a = 8'd38; b = 8'd202;  #10 
a = 8'd38; b = 8'd203;  #10 
a = 8'd38; b = 8'd204;  #10 
a = 8'd38; b = 8'd205;  #10 
a = 8'd38; b = 8'd206;  #10 
a = 8'd38; b = 8'd207;  #10 
a = 8'd38; b = 8'd208;  #10 
a = 8'd38; b = 8'd209;  #10 
a = 8'd38; b = 8'd210;  #10 
a = 8'd38; b = 8'd211;  #10 
a = 8'd38; b = 8'd212;  #10 
a = 8'd38; b = 8'd213;  #10 
a = 8'd38; b = 8'd214;  #10 
a = 8'd38; b = 8'd215;  #10 
a = 8'd38; b = 8'd216;  #10 
a = 8'd38; b = 8'd217;  #10 
a = 8'd38; b = 8'd218;  #10 
a = 8'd38; b = 8'd219;  #10 
a = 8'd38; b = 8'd220;  #10 
a = 8'd38; b = 8'd221;  #10 
a = 8'd38; b = 8'd222;  #10 
a = 8'd38; b = 8'd223;  #10 
a = 8'd38; b = 8'd224;  #10 
a = 8'd38; b = 8'd225;  #10 
a = 8'd38; b = 8'd226;  #10 
a = 8'd38; b = 8'd227;  #10 
a = 8'd38; b = 8'd228;  #10 
a = 8'd38; b = 8'd229;  #10 
a = 8'd38; b = 8'd230;  #10 
a = 8'd38; b = 8'd231;  #10 
a = 8'd38; b = 8'd232;  #10 
a = 8'd38; b = 8'd233;  #10 
a = 8'd38; b = 8'd234;  #10 
a = 8'd38; b = 8'd235;  #10 
a = 8'd38; b = 8'd236;  #10 
a = 8'd38; b = 8'd237;  #10 
a = 8'd38; b = 8'd238;  #10 
a = 8'd38; b = 8'd239;  #10 
a = 8'd38; b = 8'd240;  #10 
a = 8'd38; b = 8'd241;  #10 
a = 8'd38; b = 8'd242;  #10 
a = 8'd38; b = 8'd243;  #10 
a = 8'd38; b = 8'd244;  #10 
a = 8'd38; b = 8'd245;  #10 
a = 8'd38; b = 8'd246;  #10 
a = 8'd38; b = 8'd247;  #10 
a = 8'd38; b = 8'd248;  #10 
a = 8'd38; b = 8'd249;  #10 
a = 8'd38; b = 8'd250;  #10 
a = 8'd38; b = 8'd251;  #10 
a = 8'd38; b = 8'd252;  #10 
a = 8'd38; b = 8'd253;  #10 
a = 8'd38; b = 8'd254;  #10 
a = 8'd38; b = 8'd255;  #10 
a = 8'd39; b = 8'd0;  #10 
a = 8'd39; b = 8'd1;  #10 
a = 8'd39; b = 8'd2;  #10 
a = 8'd39; b = 8'd3;  #10 
a = 8'd39; b = 8'd4;  #10 
a = 8'd39; b = 8'd5;  #10 
a = 8'd39; b = 8'd6;  #10 
a = 8'd39; b = 8'd7;  #10 
a = 8'd39; b = 8'd8;  #10 
a = 8'd39; b = 8'd9;  #10 
a = 8'd39; b = 8'd10;  #10 
a = 8'd39; b = 8'd11;  #10 
a = 8'd39; b = 8'd12;  #10 
a = 8'd39; b = 8'd13;  #10 
a = 8'd39; b = 8'd14;  #10 
a = 8'd39; b = 8'd15;  #10 
a = 8'd39; b = 8'd16;  #10 
a = 8'd39; b = 8'd17;  #10 
a = 8'd39; b = 8'd18;  #10 
a = 8'd39; b = 8'd19;  #10 
a = 8'd39; b = 8'd20;  #10 
a = 8'd39; b = 8'd21;  #10 
a = 8'd39; b = 8'd22;  #10 
a = 8'd39; b = 8'd23;  #10 
a = 8'd39; b = 8'd24;  #10 
a = 8'd39; b = 8'd25;  #10 
a = 8'd39; b = 8'd26;  #10 
a = 8'd39; b = 8'd27;  #10 
a = 8'd39; b = 8'd28;  #10 
a = 8'd39; b = 8'd29;  #10 
a = 8'd39; b = 8'd30;  #10 
a = 8'd39; b = 8'd31;  #10 
a = 8'd39; b = 8'd32;  #10 
a = 8'd39; b = 8'd33;  #10 
a = 8'd39; b = 8'd34;  #10 
a = 8'd39; b = 8'd35;  #10 
a = 8'd39; b = 8'd36;  #10 
a = 8'd39; b = 8'd37;  #10 
a = 8'd39; b = 8'd38;  #10 
a = 8'd39; b = 8'd39;  #10 
a = 8'd39; b = 8'd40;  #10 
a = 8'd39; b = 8'd41;  #10 
a = 8'd39; b = 8'd42;  #10 
a = 8'd39; b = 8'd43;  #10 
a = 8'd39; b = 8'd44;  #10 
a = 8'd39; b = 8'd45;  #10 
a = 8'd39; b = 8'd46;  #10 
a = 8'd39; b = 8'd47;  #10 
a = 8'd39; b = 8'd48;  #10 
a = 8'd39; b = 8'd49;  #10 
a = 8'd39; b = 8'd50;  #10 
a = 8'd39; b = 8'd51;  #10 
a = 8'd39; b = 8'd52;  #10 
a = 8'd39; b = 8'd53;  #10 
a = 8'd39; b = 8'd54;  #10 
a = 8'd39; b = 8'd55;  #10 
a = 8'd39; b = 8'd56;  #10 
a = 8'd39; b = 8'd57;  #10 
a = 8'd39; b = 8'd58;  #10 
a = 8'd39; b = 8'd59;  #10 
a = 8'd39; b = 8'd60;  #10 
a = 8'd39; b = 8'd61;  #10 
a = 8'd39; b = 8'd62;  #10 
a = 8'd39; b = 8'd63;  #10 
a = 8'd39; b = 8'd64;  #10 
a = 8'd39; b = 8'd65;  #10 
a = 8'd39; b = 8'd66;  #10 
a = 8'd39; b = 8'd67;  #10 
a = 8'd39; b = 8'd68;  #10 
a = 8'd39; b = 8'd69;  #10 
a = 8'd39; b = 8'd70;  #10 
a = 8'd39; b = 8'd71;  #10 
a = 8'd39; b = 8'd72;  #10 
a = 8'd39; b = 8'd73;  #10 
a = 8'd39; b = 8'd74;  #10 
a = 8'd39; b = 8'd75;  #10 
a = 8'd39; b = 8'd76;  #10 
a = 8'd39; b = 8'd77;  #10 
a = 8'd39; b = 8'd78;  #10 
a = 8'd39; b = 8'd79;  #10 
a = 8'd39; b = 8'd80;  #10 
a = 8'd39; b = 8'd81;  #10 
a = 8'd39; b = 8'd82;  #10 
a = 8'd39; b = 8'd83;  #10 
a = 8'd39; b = 8'd84;  #10 
a = 8'd39; b = 8'd85;  #10 
a = 8'd39; b = 8'd86;  #10 
a = 8'd39; b = 8'd87;  #10 
a = 8'd39; b = 8'd88;  #10 
a = 8'd39; b = 8'd89;  #10 
a = 8'd39; b = 8'd90;  #10 
a = 8'd39; b = 8'd91;  #10 
a = 8'd39; b = 8'd92;  #10 
a = 8'd39; b = 8'd93;  #10 
a = 8'd39; b = 8'd94;  #10 
a = 8'd39; b = 8'd95;  #10 
a = 8'd39; b = 8'd96;  #10 
a = 8'd39; b = 8'd97;  #10 
a = 8'd39; b = 8'd98;  #10 
a = 8'd39; b = 8'd99;  #10 
a = 8'd39; b = 8'd100;  #10 
a = 8'd39; b = 8'd101;  #10 
a = 8'd39; b = 8'd102;  #10 
a = 8'd39; b = 8'd103;  #10 
a = 8'd39; b = 8'd104;  #10 
a = 8'd39; b = 8'd105;  #10 
a = 8'd39; b = 8'd106;  #10 
a = 8'd39; b = 8'd107;  #10 
a = 8'd39; b = 8'd108;  #10 
a = 8'd39; b = 8'd109;  #10 
a = 8'd39; b = 8'd110;  #10 
a = 8'd39; b = 8'd111;  #10 
a = 8'd39; b = 8'd112;  #10 
a = 8'd39; b = 8'd113;  #10 
a = 8'd39; b = 8'd114;  #10 
a = 8'd39; b = 8'd115;  #10 
a = 8'd39; b = 8'd116;  #10 
a = 8'd39; b = 8'd117;  #10 
a = 8'd39; b = 8'd118;  #10 
a = 8'd39; b = 8'd119;  #10 
a = 8'd39; b = 8'd120;  #10 
a = 8'd39; b = 8'd121;  #10 
a = 8'd39; b = 8'd122;  #10 
a = 8'd39; b = 8'd123;  #10 
a = 8'd39; b = 8'd124;  #10 
a = 8'd39; b = 8'd125;  #10 
a = 8'd39; b = 8'd126;  #10 
a = 8'd39; b = 8'd127;  #10 
a = 8'd39; b = 8'd128;  #10 
a = 8'd39; b = 8'd129;  #10 
a = 8'd39; b = 8'd130;  #10 
a = 8'd39; b = 8'd131;  #10 
a = 8'd39; b = 8'd132;  #10 
a = 8'd39; b = 8'd133;  #10 
a = 8'd39; b = 8'd134;  #10 
a = 8'd39; b = 8'd135;  #10 
a = 8'd39; b = 8'd136;  #10 
a = 8'd39; b = 8'd137;  #10 
a = 8'd39; b = 8'd138;  #10 
a = 8'd39; b = 8'd139;  #10 
a = 8'd39; b = 8'd140;  #10 
a = 8'd39; b = 8'd141;  #10 
a = 8'd39; b = 8'd142;  #10 
a = 8'd39; b = 8'd143;  #10 
a = 8'd39; b = 8'd144;  #10 
a = 8'd39; b = 8'd145;  #10 
a = 8'd39; b = 8'd146;  #10 
a = 8'd39; b = 8'd147;  #10 
a = 8'd39; b = 8'd148;  #10 
a = 8'd39; b = 8'd149;  #10 
a = 8'd39; b = 8'd150;  #10 
a = 8'd39; b = 8'd151;  #10 
a = 8'd39; b = 8'd152;  #10 
a = 8'd39; b = 8'd153;  #10 
a = 8'd39; b = 8'd154;  #10 
a = 8'd39; b = 8'd155;  #10 
a = 8'd39; b = 8'd156;  #10 
a = 8'd39; b = 8'd157;  #10 
a = 8'd39; b = 8'd158;  #10 
a = 8'd39; b = 8'd159;  #10 
a = 8'd39; b = 8'd160;  #10 
a = 8'd39; b = 8'd161;  #10 
a = 8'd39; b = 8'd162;  #10 
a = 8'd39; b = 8'd163;  #10 
a = 8'd39; b = 8'd164;  #10 
a = 8'd39; b = 8'd165;  #10 
a = 8'd39; b = 8'd166;  #10 
a = 8'd39; b = 8'd167;  #10 
a = 8'd39; b = 8'd168;  #10 
a = 8'd39; b = 8'd169;  #10 
a = 8'd39; b = 8'd170;  #10 
a = 8'd39; b = 8'd171;  #10 
a = 8'd39; b = 8'd172;  #10 
a = 8'd39; b = 8'd173;  #10 
a = 8'd39; b = 8'd174;  #10 
a = 8'd39; b = 8'd175;  #10 
a = 8'd39; b = 8'd176;  #10 
a = 8'd39; b = 8'd177;  #10 
a = 8'd39; b = 8'd178;  #10 
a = 8'd39; b = 8'd179;  #10 
a = 8'd39; b = 8'd180;  #10 
a = 8'd39; b = 8'd181;  #10 
a = 8'd39; b = 8'd182;  #10 
a = 8'd39; b = 8'd183;  #10 
a = 8'd39; b = 8'd184;  #10 
a = 8'd39; b = 8'd185;  #10 
a = 8'd39; b = 8'd186;  #10 
a = 8'd39; b = 8'd187;  #10 
a = 8'd39; b = 8'd188;  #10 
a = 8'd39; b = 8'd189;  #10 
a = 8'd39; b = 8'd190;  #10 
a = 8'd39; b = 8'd191;  #10 
a = 8'd39; b = 8'd192;  #10 
a = 8'd39; b = 8'd193;  #10 
a = 8'd39; b = 8'd194;  #10 
a = 8'd39; b = 8'd195;  #10 
a = 8'd39; b = 8'd196;  #10 
a = 8'd39; b = 8'd197;  #10 
a = 8'd39; b = 8'd198;  #10 
a = 8'd39; b = 8'd199;  #10 
a = 8'd39; b = 8'd200;  #10 
a = 8'd39; b = 8'd201;  #10 
a = 8'd39; b = 8'd202;  #10 
a = 8'd39; b = 8'd203;  #10 
a = 8'd39; b = 8'd204;  #10 
a = 8'd39; b = 8'd205;  #10 
a = 8'd39; b = 8'd206;  #10 
a = 8'd39; b = 8'd207;  #10 
a = 8'd39; b = 8'd208;  #10 
a = 8'd39; b = 8'd209;  #10 
a = 8'd39; b = 8'd210;  #10 
a = 8'd39; b = 8'd211;  #10 
a = 8'd39; b = 8'd212;  #10 
a = 8'd39; b = 8'd213;  #10 
a = 8'd39; b = 8'd214;  #10 
a = 8'd39; b = 8'd215;  #10 
a = 8'd39; b = 8'd216;  #10 
a = 8'd39; b = 8'd217;  #10 
a = 8'd39; b = 8'd218;  #10 
a = 8'd39; b = 8'd219;  #10 
a = 8'd39; b = 8'd220;  #10 
a = 8'd39; b = 8'd221;  #10 
a = 8'd39; b = 8'd222;  #10 
a = 8'd39; b = 8'd223;  #10 
a = 8'd39; b = 8'd224;  #10 
a = 8'd39; b = 8'd225;  #10 
a = 8'd39; b = 8'd226;  #10 
a = 8'd39; b = 8'd227;  #10 
a = 8'd39; b = 8'd228;  #10 
a = 8'd39; b = 8'd229;  #10 
a = 8'd39; b = 8'd230;  #10 
a = 8'd39; b = 8'd231;  #10 
a = 8'd39; b = 8'd232;  #10 
a = 8'd39; b = 8'd233;  #10 
a = 8'd39; b = 8'd234;  #10 
a = 8'd39; b = 8'd235;  #10 
a = 8'd39; b = 8'd236;  #10 
a = 8'd39; b = 8'd237;  #10 
a = 8'd39; b = 8'd238;  #10 
a = 8'd39; b = 8'd239;  #10 
a = 8'd39; b = 8'd240;  #10 
a = 8'd39; b = 8'd241;  #10 
a = 8'd39; b = 8'd242;  #10 
a = 8'd39; b = 8'd243;  #10 
a = 8'd39; b = 8'd244;  #10 
a = 8'd39; b = 8'd245;  #10 
a = 8'd39; b = 8'd246;  #10 
a = 8'd39; b = 8'd247;  #10 
a = 8'd39; b = 8'd248;  #10 
a = 8'd39; b = 8'd249;  #10 
a = 8'd39; b = 8'd250;  #10 
a = 8'd39; b = 8'd251;  #10 
a = 8'd39; b = 8'd252;  #10 
a = 8'd39; b = 8'd253;  #10 
a = 8'd39; b = 8'd254;  #10 
a = 8'd39; b = 8'd255;  #10 
a = 8'd40; b = 8'd0;  #10 
a = 8'd40; b = 8'd1;  #10 
a = 8'd40; b = 8'd2;  #10 
a = 8'd40; b = 8'd3;  #10 
a = 8'd40; b = 8'd4;  #10 
a = 8'd40; b = 8'd5;  #10 
a = 8'd40; b = 8'd6;  #10 
a = 8'd40; b = 8'd7;  #10 
a = 8'd40; b = 8'd8;  #10 
a = 8'd40; b = 8'd9;  #10 
a = 8'd40; b = 8'd10;  #10 
a = 8'd40; b = 8'd11;  #10 
a = 8'd40; b = 8'd12;  #10 
a = 8'd40; b = 8'd13;  #10 
a = 8'd40; b = 8'd14;  #10 
a = 8'd40; b = 8'd15;  #10 
a = 8'd40; b = 8'd16;  #10 
a = 8'd40; b = 8'd17;  #10 
a = 8'd40; b = 8'd18;  #10 
a = 8'd40; b = 8'd19;  #10 
a = 8'd40; b = 8'd20;  #10 
a = 8'd40; b = 8'd21;  #10 
a = 8'd40; b = 8'd22;  #10 
a = 8'd40; b = 8'd23;  #10 
a = 8'd40; b = 8'd24;  #10 
a = 8'd40; b = 8'd25;  #10 
a = 8'd40; b = 8'd26;  #10 
a = 8'd40; b = 8'd27;  #10 
a = 8'd40; b = 8'd28;  #10 
a = 8'd40; b = 8'd29;  #10 
a = 8'd40; b = 8'd30;  #10 
a = 8'd40; b = 8'd31;  #10 
a = 8'd40; b = 8'd32;  #10 
a = 8'd40; b = 8'd33;  #10 
a = 8'd40; b = 8'd34;  #10 
a = 8'd40; b = 8'd35;  #10 
a = 8'd40; b = 8'd36;  #10 
a = 8'd40; b = 8'd37;  #10 
a = 8'd40; b = 8'd38;  #10 
a = 8'd40; b = 8'd39;  #10 
a = 8'd40; b = 8'd40;  #10 
a = 8'd40; b = 8'd41;  #10 
a = 8'd40; b = 8'd42;  #10 
a = 8'd40; b = 8'd43;  #10 
a = 8'd40; b = 8'd44;  #10 
a = 8'd40; b = 8'd45;  #10 
a = 8'd40; b = 8'd46;  #10 
a = 8'd40; b = 8'd47;  #10 
a = 8'd40; b = 8'd48;  #10 
a = 8'd40; b = 8'd49;  #10 
a = 8'd40; b = 8'd50;  #10 
a = 8'd40; b = 8'd51;  #10 
a = 8'd40; b = 8'd52;  #10 
a = 8'd40; b = 8'd53;  #10 
a = 8'd40; b = 8'd54;  #10 
a = 8'd40; b = 8'd55;  #10 
a = 8'd40; b = 8'd56;  #10 
a = 8'd40; b = 8'd57;  #10 
a = 8'd40; b = 8'd58;  #10 
a = 8'd40; b = 8'd59;  #10 
a = 8'd40; b = 8'd60;  #10 
a = 8'd40; b = 8'd61;  #10 
a = 8'd40; b = 8'd62;  #10 
a = 8'd40; b = 8'd63;  #10 
a = 8'd40; b = 8'd64;  #10 
a = 8'd40; b = 8'd65;  #10 
a = 8'd40; b = 8'd66;  #10 
a = 8'd40; b = 8'd67;  #10 
a = 8'd40; b = 8'd68;  #10 
a = 8'd40; b = 8'd69;  #10 
a = 8'd40; b = 8'd70;  #10 
a = 8'd40; b = 8'd71;  #10 
a = 8'd40; b = 8'd72;  #10 
a = 8'd40; b = 8'd73;  #10 
a = 8'd40; b = 8'd74;  #10 
a = 8'd40; b = 8'd75;  #10 
a = 8'd40; b = 8'd76;  #10 
a = 8'd40; b = 8'd77;  #10 
a = 8'd40; b = 8'd78;  #10 
a = 8'd40; b = 8'd79;  #10 
a = 8'd40; b = 8'd80;  #10 
a = 8'd40; b = 8'd81;  #10 
a = 8'd40; b = 8'd82;  #10 
a = 8'd40; b = 8'd83;  #10 
a = 8'd40; b = 8'd84;  #10 
a = 8'd40; b = 8'd85;  #10 
a = 8'd40; b = 8'd86;  #10 
a = 8'd40; b = 8'd87;  #10 
a = 8'd40; b = 8'd88;  #10 
a = 8'd40; b = 8'd89;  #10 
a = 8'd40; b = 8'd90;  #10 
a = 8'd40; b = 8'd91;  #10 
a = 8'd40; b = 8'd92;  #10 
a = 8'd40; b = 8'd93;  #10 
a = 8'd40; b = 8'd94;  #10 
a = 8'd40; b = 8'd95;  #10 
a = 8'd40; b = 8'd96;  #10 
a = 8'd40; b = 8'd97;  #10 
a = 8'd40; b = 8'd98;  #10 
a = 8'd40; b = 8'd99;  #10 
a = 8'd40; b = 8'd100;  #10 
a = 8'd40; b = 8'd101;  #10 
a = 8'd40; b = 8'd102;  #10 
a = 8'd40; b = 8'd103;  #10 
a = 8'd40; b = 8'd104;  #10 
a = 8'd40; b = 8'd105;  #10 
a = 8'd40; b = 8'd106;  #10 
a = 8'd40; b = 8'd107;  #10 
a = 8'd40; b = 8'd108;  #10 
a = 8'd40; b = 8'd109;  #10 
a = 8'd40; b = 8'd110;  #10 
a = 8'd40; b = 8'd111;  #10 
a = 8'd40; b = 8'd112;  #10 
a = 8'd40; b = 8'd113;  #10 
a = 8'd40; b = 8'd114;  #10 
a = 8'd40; b = 8'd115;  #10 
a = 8'd40; b = 8'd116;  #10 
a = 8'd40; b = 8'd117;  #10 
a = 8'd40; b = 8'd118;  #10 
a = 8'd40; b = 8'd119;  #10 
a = 8'd40; b = 8'd120;  #10 
a = 8'd40; b = 8'd121;  #10 
a = 8'd40; b = 8'd122;  #10 
a = 8'd40; b = 8'd123;  #10 
a = 8'd40; b = 8'd124;  #10 
a = 8'd40; b = 8'd125;  #10 
a = 8'd40; b = 8'd126;  #10 
a = 8'd40; b = 8'd127;  #10 
a = 8'd40; b = 8'd128;  #10 
a = 8'd40; b = 8'd129;  #10 
a = 8'd40; b = 8'd130;  #10 
a = 8'd40; b = 8'd131;  #10 
a = 8'd40; b = 8'd132;  #10 
a = 8'd40; b = 8'd133;  #10 
a = 8'd40; b = 8'd134;  #10 
a = 8'd40; b = 8'd135;  #10 
a = 8'd40; b = 8'd136;  #10 
a = 8'd40; b = 8'd137;  #10 
a = 8'd40; b = 8'd138;  #10 
a = 8'd40; b = 8'd139;  #10 
a = 8'd40; b = 8'd140;  #10 
a = 8'd40; b = 8'd141;  #10 
a = 8'd40; b = 8'd142;  #10 
a = 8'd40; b = 8'd143;  #10 
a = 8'd40; b = 8'd144;  #10 
a = 8'd40; b = 8'd145;  #10 
a = 8'd40; b = 8'd146;  #10 
a = 8'd40; b = 8'd147;  #10 
a = 8'd40; b = 8'd148;  #10 
a = 8'd40; b = 8'd149;  #10 
a = 8'd40; b = 8'd150;  #10 
a = 8'd40; b = 8'd151;  #10 
a = 8'd40; b = 8'd152;  #10 
a = 8'd40; b = 8'd153;  #10 
a = 8'd40; b = 8'd154;  #10 
a = 8'd40; b = 8'd155;  #10 
a = 8'd40; b = 8'd156;  #10 
a = 8'd40; b = 8'd157;  #10 
a = 8'd40; b = 8'd158;  #10 
a = 8'd40; b = 8'd159;  #10 
a = 8'd40; b = 8'd160;  #10 
a = 8'd40; b = 8'd161;  #10 
a = 8'd40; b = 8'd162;  #10 
a = 8'd40; b = 8'd163;  #10 
a = 8'd40; b = 8'd164;  #10 
a = 8'd40; b = 8'd165;  #10 
a = 8'd40; b = 8'd166;  #10 
a = 8'd40; b = 8'd167;  #10 
a = 8'd40; b = 8'd168;  #10 
a = 8'd40; b = 8'd169;  #10 
a = 8'd40; b = 8'd170;  #10 
a = 8'd40; b = 8'd171;  #10 
a = 8'd40; b = 8'd172;  #10 
a = 8'd40; b = 8'd173;  #10 
a = 8'd40; b = 8'd174;  #10 
a = 8'd40; b = 8'd175;  #10 
a = 8'd40; b = 8'd176;  #10 
a = 8'd40; b = 8'd177;  #10 
a = 8'd40; b = 8'd178;  #10 
a = 8'd40; b = 8'd179;  #10 
a = 8'd40; b = 8'd180;  #10 
a = 8'd40; b = 8'd181;  #10 
a = 8'd40; b = 8'd182;  #10 
a = 8'd40; b = 8'd183;  #10 
a = 8'd40; b = 8'd184;  #10 
a = 8'd40; b = 8'd185;  #10 
a = 8'd40; b = 8'd186;  #10 
a = 8'd40; b = 8'd187;  #10 
a = 8'd40; b = 8'd188;  #10 
a = 8'd40; b = 8'd189;  #10 
a = 8'd40; b = 8'd190;  #10 
a = 8'd40; b = 8'd191;  #10 
a = 8'd40; b = 8'd192;  #10 
a = 8'd40; b = 8'd193;  #10 
a = 8'd40; b = 8'd194;  #10 
a = 8'd40; b = 8'd195;  #10 
a = 8'd40; b = 8'd196;  #10 
a = 8'd40; b = 8'd197;  #10 
a = 8'd40; b = 8'd198;  #10 
a = 8'd40; b = 8'd199;  #10 
a = 8'd40; b = 8'd200;  #10 
a = 8'd40; b = 8'd201;  #10 
a = 8'd40; b = 8'd202;  #10 
a = 8'd40; b = 8'd203;  #10 
a = 8'd40; b = 8'd204;  #10 
a = 8'd40; b = 8'd205;  #10 
a = 8'd40; b = 8'd206;  #10 
a = 8'd40; b = 8'd207;  #10 
a = 8'd40; b = 8'd208;  #10 
a = 8'd40; b = 8'd209;  #10 
a = 8'd40; b = 8'd210;  #10 
a = 8'd40; b = 8'd211;  #10 
a = 8'd40; b = 8'd212;  #10 
a = 8'd40; b = 8'd213;  #10 
a = 8'd40; b = 8'd214;  #10 
a = 8'd40; b = 8'd215;  #10 
a = 8'd40; b = 8'd216;  #10 
a = 8'd40; b = 8'd217;  #10 
a = 8'd40; b = 8'd218;  #10 
a = 8'd40; b = 8'd219;  #10 
a = 8'd40; b = 8'd220;  #10 
a = 8'd40; b = 8'd221;  #10 
a = 8'd40; b = 8'd222;  #10 
a = 8'd40; b = 8'd223;  #10 
a = 8'd40; b = 8'd224;  #10 
a = 8'd40; b = 8'd225;  #10 
a = 8'd40; b = 8'd226;  #10 
a = 8'd40; b = 8'd227;  #10 
a = 8'd40; b = 8'd228;  #10 
a = 8'd40; b = 8'd229;  #10 
a = 8'd40; b = 8'd230;  #10 
a = 8'd40; b = 8'd231;  #10 
a = 8'd40; b = 8'd232;  #10 
a = 8'd40; b = 8'd233;  #10 
a = 8'd40; b = 8'd234;  #10 
a = 8'd40; b = 8'd235;  #10 
a = 8'd40; b = 8'd236;  #10 
a = 8'd40; b = 8'd237;  #10 
a = 8'd40; b = 8'd238;  #10 
a = 8'd40; b = 8'd239;  #10 
a = 8'd40; b = 8'd240;  #10 
a = 8'd40; b = 8'd241;  #10 
a = 8'd40; b = 8'd242;  #10 
a = 8'd40; b = 8'd243;  #10 
a = 8'd40; b = 8'd244;  #10 
a = 8'd40; b = 8'd245;  #10 
a = 8'd40; b = 8'd246;  #10 
a = 8'd40; b = 8'd247;  #10 
a = 8'd40; b = 8'd248;  #10 
a = 8'd40; b = 8'd249;  #10 
a = 8'd40; b = 8'd250;  #10 
a = 8'd40; b = 8'd251;  #10 
a = 8'd40; b = 8'd252;  #10 
a = 8'd40; b = 8'd253;  #10 
a = 8'd40; b = 8'd254;  #10 
a = 8'd40; b = 8'd255;  #10 
a = 8'd41; b = 8'd0;  #10 
a = 8'd41; b = 8'd1;  #10 
a = 8'd41; b = 8'd2;  #10 
a = 8'd41; b = 8'd3;  #10 
a = 8'd41; b = 8'd4;  #10 
a = 8'd41; b = 8'd5;  #10 
a = 8'd41; b = 8'd6;  #10 
a = 8'd41; b = 8'd7;  #10 
a = 8'd41; b = 8'd8;  #10 
a = 8'd41; b = 8'd9;  #10 
a = 8'd41; b = 8'd10;  #10 
a = 8'd41; b = 8'd11;  #10 
a = 8'd41; b = 8'd12;  #10 
a = 8'd41; b = 8'd13;  #10 
a = 8'd41; b = 8'd14;  #10 
a = 8'd41; b = 8'd15;  #10 
a = 8'd41; b = 8'd16;  #10 
a = 8'd41; b = 8'd17;  #10 
a = 8'd41; b = 8'd18;  #10 
a = 8'd41; b = 8'd19;  #10 
a = 8'd41; b = 8'd20;  #10 
a = 8'd41; b = 8'd21;  #10 
a = 8'd41; b = 8'd22;  #10 
a = 8'd41; b = 8'd23;  #10 
a = 8'd41; b = 8'd24;  #10 
a = 8'd41; b = 8'd25;  #10 
a = 8'd41; b = 8'd26;  #10 
a = 8'd41; b = 8'd27;  #10 
a = 8'd41; b = 8'd28;  #10 
a = 8'd41; b = 8'd29;  #10 
a = 8'd41; b = 8'd30;  #10 
a = 8'd41; b = 8'd31;  #10 
a = 8'd41; b = 8'd32;  #10 
a = 8'd41; b = 8'd33;  #10 
a = 8'd41; b = 8'd34;  #10 
a = 8'd41; b = 8'd35;  #10 
a = 8'd41; b = 8'd36;  #10 
a = 8'd41; b = 8'd37;  #10 
a = 8'd41; b = 8'd38;  #10 
a = 8'd41; b = 8'd39;  #10 
a = 8'd41; b = 8'd40;  #10 
a = 8'd41; b = 8'd41;  #10 
a = 8'd41; b = 8'd42;  #10 
a = 8'd41; b = 8'd43;  #10 
a = 8'd41; b = 8'd44;  #10 
a = 8'd41; b = 8'd45;  #10 
a = 8'd41; b = 8'd46;  #10 
a = 8'd41; b = 8'd47;  #10 
a = 8'd41; b = 8'd48;  #10 
a = 8'd41; b = 8'd49;  #10 
a = 8'd41; b = 8'd50;  #10 
a = 8'd41; b = 8'd51;  #10 
a = 8'd41; b = 8'd52;  #10 
a = 8'd41; b = 8'd53;  #10 
a = 8'd41; b = 8'd54;  #10 
a = 8'd41; b = 8'd55;  #10 
a = 8'd41; b = 8'd56;  #10 
a = 8'd41; b = 8'd57;  #10 
a = 8'd41; b = 8'd58;  #10 
a = 8'd41; b = 8'd59;  #10 
a = 8'd41; b = 8'd60;  #10 
a = 8'd41; b = 8'd61;  #10 
a = 8'd41; b = 8'd62;  #10 
a = 8'd41; b = 8'd63;  #10 
a = 8'd41; b = 8'd64;  #10 
a = 8'd41; b = 8'd65;  #10 
a = 8'd41; b = 8'd66;  #10 
a = 8'd41; b = 8'd67;  #10 
a = 8'd41; b = 8'd68;  #10 
a = 8'd41; b = 8'd69;  #10 
a = 8'd41; b = 8'd70;  #10 
a = 8'd41; b = 8'd71;  #10 
a = 8'd41; b = 8'd72;  #10 
a = 8'd41; b = 8'd73;  #10 
a = 8'd41; b = 8'd74;  #10 
a = 8'd41; b = 8'd75;  #10 
a = 8'd41; b = 8'd76;  #10 
a = 8'd41; b = 8'd77;  #10 
a = 8'd41; b = 8'd78;  #10 
a = 8'd41; b = 8'd79;  #10 
a = 8'd41; b = 8'd80;  #10 
a = 8'd41; b = 8'd81;  #10 
a = 8'd41; b = 8'd82;  #10 
a = 8'd41; b = 8'd83;  #10 
a = 8'd41; b = 8'd84;  #10 
a = 8'd41; b = 8'd85;  #10 
a = 8'd41; b = 8'd86;  #10 
a = 8'd41; b = 8'd87;  #10 
a = 8'd41; b = 8'd88;  #10 
a = 8'd41; b = 8'd89;  #10 
a = 8'd41; b = 8'd90;  #10 
a = 8'd41; b = 8'd91;  #10 
a = 8'd41; b = 8'd92;  #10 
a = 8'd41; b = 8'd93;  #10 
a = 8'd41; b = 8'd94;  #10 
a = 8'd41; b = 8'd95;  #10 
a = 8'd41; b = 8'd96;  #10 
a = 8'd41; b = 8'd97;  #10 
a = 8'd41; b = 8'd98;  #10 
a = 8'd41; b = 8'd99;  #10 
a = 8'd41; b = 8'd100;  #10 
a = 8'd41; b = 8'd101;  #10 
a = 8'd41; b = 8'd102;  #10 
a = 8'd41; b = 8'd103;  #10 
a = 8'd41; b = 8'd104;  #10 
a = 8'd41; b = 8'd105;  #10 
a = 8'd41; b = 8'd106;  #10 
a = 8'd41; b = 8'd107;  #10 
a = 8'd41; b = 8'd108;  #10 
a = 8'd41; b = 8'd109;  #10 
a = 8'd41; b = 8'd110;  #10 
a = 8'd41; b = 8'd111;  #10 
a = 8'd41; b = 8'd112;  #10 
a = 8'd41; b = 8'd113;  #10 
a = 8'd41; b = 8'd114;  #10 
a = 8'd41; b = 8'd115;  #10 
a = 8'd41; b = 8'd116;  #10 
a = 8'd41; b = 8'd117;  #10 
a = 8'd41; b = 8'd118;  #10 
a = 8'd41; b = 8'd119;  #10 
a = 8'd41; b = 8'd120;  #10 
a = 8'd41; b = 8'd121;  #10 
a = 8'd41; b = 8'd122;  #10 
a = 8'd41; b = 8'd123;  #10 
a = 8'd41; b = 8'd124;  #10 
a = 8'd41; b = 8'd125;  #10 
a = 8'd41; b = 8'd126;  #10 
a = 8'd41; b = 8'd127;  #10 
a = 8'd41; b = 8'd128;  #10 
a = 8'd41; b = 8'd129;  #10 
a = 8'd41; b = 8'd130;  #10 
a = 8'd41; b = 8'd131;  #10 
a = 8'd41; b = 8'd132;  #10 
a = 8'd41; b = 8'd133;  #10 
a = 8'd41; b = 8'd134;  #10 
a = 8'd41; b = 8'd135;  #10 
a = 8'd41; b = 8'd136;  #10 
a = 8'd41; b = 8'd137;  #10 
a = 8'd41; b = 8'd138;  #10 
a = 8'd41; b = 8'd139;  #10 
a = 8'd41; b = 8'd140;  #10 
a = 8'd41; b = 8'd141;  #10 
a = 8'd41; b = 8'd142;  #10 
a = 8'd41; b = 8'd143;  #10 
a = 8'd41; b = 8'd144;  #10 
a = 8'd41; b = 8'd145;  #10 
a = 8'd41; b = 8'd146;  #10 
a = 8'd41; b = 8'd147;  #10 
a = 8'd41; b = 8'd148;  #10 
a = 8'd41; b = 8'd149;  #10 
a = 8'd41; b = 8'd150;  #10 
a = 8'd41; b = 8'd151;  #10 
a = 8'd41; b = 8'd152;  #10 
a = 8'd41; b = 8'd153;  #10 
a = 8'd41; b = 8'd154;  #10 
a = 8'd41; b = 8'd155;  #10 
a = 8'd41; b = 8'd156;  #10 
a = 8'd41; b = 8'd157;  #10 
a = 8'd41; b = 8'd158;  #10 
a = 8'd41; b = 8'd159;  #10 
a = 8'd41; b = 8'd160;  #10 
a = 8'd41; b = 8'd161;  #10 
a = 8'd41; b = 8'd162;  #10 
a = 8'd41; b = 8'd163;  #10 
a = 8'd41; b = 8'd164;  #10 
a = 8'd41; b = 8'd165;  #10 
a = 8'd41; b = 8'd166;  #10 
a = 8'd41; b = 8'd167;  #10 
a = 8'd41; b = 8'd168;  #10 
a = 8'd41; b = 8'd169;  #10 
a = 8'd41; b = 8'd170;  #10 
a = 8'd41; b = 8'd171;  #10 
a = 8'd41; b = 8'd172;  #10 
a = 8'd41; b = 8'd173;  #10 
a = 8'd41; b = 8'd174;  #10 
a = 8'd41; b = 8'd175;  #10 
a = 8'd41; b = 8'd176;  #10 
a = 8'd41; b = 8'd177;  #10 
a = 8'd41; b = 8'd178;  #10 
a = 8'd41; b = 8'd179;  #10 
a = 8'd41; b = 8'd180;  #10 
a = 8'd41; b = 8'd181;  #10 
a = 8'd41; b = 8'd182;  #10 
a = 8'd41; b = 8'd183;  #10 
a = 8'd41; b = 8'd184;  #10 
a = 8'd41; b = 8'd185;  #10 
a = 8'd41; b = 8'd186;  #10 
a = 8'd41; b = 8'd187;  #10 
a = 8'd41; b = 8'd188;  #10 
a = 8'd41; b = 8'd189;  #10 
a = 8'd41; b = 8'd190;  #10 
a = 8'd41; b = 8'd191;  #10 
a = 8'd41; b = 8'd192;  #10 
a = 8'd41; b = 8'd193;  #10 
a = 8'd41; b = 8'd194;  #10 
a = 8'd41; b = 8'd195;  #10 
a = 8'd41; b = 8'd196;  #10 
a = 8'd41; b = 8'd197;  #10 
a = 8'd41; b = 8'd198;  #10 
a = 8'd41; b = 8'd199;  #10 
a = 8'd41; b = 8'd200;  #10 
a = 8'd41; b = 8'd201;  #10 
a = 8'd41; b = 8'd202;  #10 
a = 8'd41; b = 8'd203;  #10 
a = 8'd41; b = 8'd204;  #10 
a = 8'd41; b = 8'd205;  #10 
a = 8'd41; b = 8'd206;  #10 
a = 8'd41; b = 8'd207;  #10 
a = 8'd41; b = 8'd208;  #10 
a = 8'd41; b = 8'd209;  #10 
a = 8'd41; b = 8'd210;  #10 
a = 8'd41; b = 8'd211;  #10 
a = 8'd41; b = 8'd212;  #10 
a = 8'd41; b = 8'd213;  #10 
a = 8'd41; b = 8'd214;  #10 
a = 8'd41; b = 8'd215;  #10 
a = 8'd41; b = 8'd216;  #10 
a = 8'd41; b = 8'd217;  #10 
a = 8'd41; b = 8'd218;  #10 
a = 8'd41; b = 8'd219;  #10 
a = 8'd41; b = 8'd220;  #10 
a = 8'd41; b = 8'd221;  #10 
a = 8'd41; b = 8'd222;  #10 
a = 8'd41; b = 8'd223;  #10 
a = 8'd41; b = 8'd224;  #10 
a = 8'd41; b = 8'd225;  #10 
a = 8'd41; b = 8'd226;  #10 
a = 8'd41; b = 8'd227;  #10 
a = 8'd41; b = 8'd228;  #10 
a = 8'd41; b = 8'd229;  #10 
a = 8'd41; b = 8'd230;  #10 
a = 8'd41; b = 8'd231;  #10 
a = 8'd41; b = 8'd232;  #10 
a = 8'd41; b = 8'd233;  #10 
a = 8'd41; b = 8'd234;  #10 
a = 8'd41; b = 8'd235;  #10 
a = 8'd41; b = 8'd236;  #10 
a = 8'd41; b = 8'd237;  #10 
a = 8'd41; b = 8'd238;  #10 
a = 8'd41; b = 8'd239;  #10 
a = 8'd41; b = 8'd240;  #10 
a = 8'd41; b = 8'd241;  #10 
a = 8'd41; b = 8'd242;  #10 
a = 8'd41; b = 8'd243;  #10 
a = 8'd41; b = 8'd244;  #10 
a = 8'd41; b = 8'd245;  #10 
a = 8'd41; b = 8'd246;  #10 
a = 8'd41; b = 8'd247;  #10 
a = 8'd41; b = 8'd248;  #10 
a = 8'd41; b = 8'd249;  #10 
a = 8'd41; b = 8'd250;  #10 
a = 8'd41; b = 8'd251;  #10 
a = 8'd41; b = 8'd252;  #10 
a = 8'd41; b = 8'd253;  #10 
a = 8'd41; b = 8'd254;  #10 
a = 8'd41; b = 8'd255;  #10 
a = 8'd42; b = 8'd0;  #10 
a = 8'd42; b = 8'd1;  #10 
a = 8'd42; b = 8'd2;  #10 
a = 8'd42; b = 8'd3;  #10 
a = 8'd42; b = 8'd4;  #10 
a = 8'd42; b = 8'd5;  #10 
a = 8'd42; b = 8'd6;  #10 
a = 8'd42; b = 8'd7;  #10 
a = 8'd42; b = 8'd8;  #10 
a = 8'd42; b = 8'd9;  #10 
a = 8'd42; b = 8'd10;  #10 
a = 8'd42; b = 8'd11;  #10 
a = 8'd42; b = 8'd12;  #10 
a = 8'd42; b = 8'd13;  #10 
a = 8'd42; b = 8'd14;  #10 
a = 8'd42; b = 8'd15;  #10 
a = 8'd42; b = 8'd16;  #10 
a = 8'd42; b = 8'd17;  #10 
a = 8'd42; b = 8'd18;  #10 
a = 8'd42; b = 8'd19;  #10 
a = 8'd42; b = 8'd20;  #10 
a = 8'd42; b = 8'd21;  #10 
a = 8'd42; b = 8'd22;  #10 
a = 8'd42; b = 8'd23;  #10 
a = 8'd42; b = 8'd24;  #10 
a = 8'd42; b = 8'd25;  #10 
a = 8'd42; b = 8'd26;  #10 
a = 8'd42; b = 8'd27;  #10 
a = 8'd42; b = 8'd28;  #10 
a = 8'd42; b = 8'd29;  #10 
a = 8'd42; b = 8'd30;  #10 
a = 8'd42; b = 8'd31;  #10 
a = 8'd42; b = 8'd32;  #10 
a = 8'd42; b = 8'd33;  #10 
a = 8'd42; b = 8'd34;  #10 
a = 8'd42; b = 8'd35;  #10 
a = 8'd42; b = 8'd36;  #10 
a = 8'd42; b = 8'd37;  #10 
a = 8'd42; b = 8'd38;  #10 
a = 8'd42; b = 8'd39;  #10 
a = 8'd42; b = 8'd40;  #10 
a = 8'd42; b = 8'd41;  #10 
a = 8'd42; b = 8'd42;  #10 
a = 8'd42; b = 8'd43;  #10 
a = 8'd42; b = 8'd44;  #10 
a = 8'd42; b = 8'd45;  #10 
a = 8'd42; b = 8'd46;  #10 
a = 8'd42; b = 8'd47;  #10 
a = 8'd42; b = 8'd48;  #10 
a = 8'd42; b = 8'd49;  #10 
a = 8'd42; b = 8'd50;  #10 
a = 8'd42; b = 8'd51;  #10 
a = 8'd42; b = 8'd52;  #10 
a = 8'd42; b = 8'd53;  #10 
a = 8'd42; b = 8'd54;  #10 
a = 8'd42; b = 8'd55;  #10 
a = 8'd42; b = 8'd56;  #10 
a = 8'd42; b = 8'd57;  #10 
a = 8'd42; b = 8'd58;  #10 
a = 8'd42; b = 8'd59;  #10 
a = 8'd42; b = 8'd60;  #10 
a = 8'd42; b = 8'd61;  #10 
a = 8'd42; b = 8'd62;  #10 
a = 8'd42; b = 8'd63;  #10 
a = 8'd42; b = 8'd64;  #10 
a = 8'd42; b = 8'd65;  #10 
a = 8'd42; b = 8'd66;  #10 
a = 8'd42; b = 8'd67;  #10 
a = 8'd42; b = 8'd68;  #10 
a = 8'd42; b = 8'd69;  #10 
a = 8'd42; b = 8'd70;  #10 
a = 8'd42; b = 8'd71;  #10 
a = 8'd42; b = 8'd72;  #10 
a = 8'd42; b = 8'd73;  #10 
a = 8'd42; b = 8'd74;  #10 
a = 8'd42; b = 8'd75;  #10 
a = 8'd42; b = 8'd76;  #10 
a = 8'd42; b = 8'd77;  #10 
a = 8'd42; b = 8'd78;  #10 
a = 8'd42; b = 8'd79;  #10 
a = 8'd42; b = 8'd80;  #10 
a = 8'd42; b = 8'd81;  #10 
a = 8'd42; b = 8'd82;  #10 
a = 8'd42; b = 8'd83;  #10 
a = 8'd42; b = 8'd84;  #10 
a = 8'd42; b = 8'd85;  #10 
a = 8'd42; b = 8'd86;  #10 
a = 8'd42; b = 8'd87;  #10 
a = 8'd42; b = 8'd88;  #10 
a = 8'd42; b = 8'd89;  #10 
a = 8'd42; b = 8'd90;  #10 
a = 8'd42; b = 8'd91;  #10 
a = 8'd42; b = 8'd92;  #10 
a = 8'd42; b = 8'd93;  #10 
a = 8'd42; b = 8'd94;  #10 
a = 8'd42; b = 8'd95;  #10 
a = 8'd42; b = 8'd96;  #10 
a = 8'd42; b = 8'd97;  #10 
a = 8'd42; b = 8'd98;  #10 
a = 8'd42; b = 8'd99;  #10 
a = 8'd42; b = 8'd100;  #10 
a = 8'd42; b = 8'd101;  #10 
a = 8'd42; b = 8'd102;  #10 
a = 8'd42; b = 8'd103;  #10 
a = 8'd42; b = 8'd104;  #10 
a = 8'd42; b = 8'd105;  #10 
a = 8'd42; b = 8'd106;  #10 
a = 8'd42; b = 8'd107;  #10 
a = 8'd42; b = 8'd108;  #10 
a = 8'd42; b = 8'd109;  #10 
a = 8'd42; b = 8'd110;  #10 
a = 8'd42; b = 8'd111;  #10 
a = 8'd42; b = 8'd112;  #10 
a = 8'd42; b = 8'd113;  #10 
a = 8'd42; b = 8'd114;  #10 
a = 8'd42; b = 8'd115;  #10 
a = 8'd42; b = 8'd116;  #10 
a = 8'd42; b = 8'd117;  #10 
a = 8'd42; b = 8'd118;  #10 
a = 8'd42; b = 8'd119;  #10 
a = 8'd42; b = 8'd120;  #10 
a = 8'd42; b = 8'd121;  #10 
a = 8'd42; b = 8'd122;  #10 
a = 8'd42; b = 8'd123;  #10 
a = 8'd42; b = 8'd124;  #10 
a = 8'd42; b = 8'd125;  #10 
a = 8'd42; b = 8'd126;  #10 
a = 8'd42; b = 8'd127;  #10 
a = 8'd42; b = 8'd128;  #10 
a = 8'd42; b = 8'd129;  #10 
a = 8'd42; b = 8'd130;  #10 
a = 8'd42; b = 8'd131;  #10 
a = 8'd42; b = 8'd132;  #10 
a = 8'd42; b = 8'd133;  #10 
a = 8'd42; b = 8'd134;  #10 
a = 8'd42; b = 8'd135;  #10 
a = 8'd42; b = 8'd136;  #10 
a = 8'd42; b = 8'd137;  #10 
a = 8'd42; b = 8'd138;  #10 
a = 8'd42; b = 8'd139;  #10 
a = 8'd42; b = 8'd140;  #10 
a = 8'd42; b = 8'd141;  #10 
a = 8'd42; b = 8'd142;  #10 
a = 8'd42; b = 8'd143;  #10 
a = 8'd42; b = 8'd144;  #10 
a = 8'd42; b = 8'd145;  #10 
a = 8'd42; b = 8'd146;  #10 
a = 8'd42; b = 8'd147;  #10 
a = 8'd42; b = 8'd148;  #10 
a = 8'd42; b = 8'd149;  #10 
a = 8'd42; b = 8'd150;  #10 
a = 8'd42; b = 8'd151;  #10 
a = 8'd42; b = 8'd152;  #10 
a = 8'd42; b = 8'd153;  #10 
a = 8'd42; b = 8'd154;  #10 
a = 8'd42; b = 8'd155;  #10 
a = 8'd42; b = 8'd156;  #10 
a = 8'd42; b = 8'd157;  #10 
a = 8'd42; b = 8'd158;  #10 
a = 8'd42; b = 8'd159;  #10 
a = 8'd42; b = 8'd160;  #10 
a = 8'd42; b = 8'd161;  #10 
a = 8'd42; b = 8'd162;  #10 
a = 8'd42; b = 8'd163;  #10 
a = 8'd42; b = 8'd164;  #10 
a = 8'd42; b = 8'd165;  #10 
a = 8'd42; b = 8'd166;  #10 
a = 8'd42; b = 8'd167;  #10 
a = 8'd42; b = 8'd168;  #10 
a = 8'd42; b = 8'd169;  #10 
a = 8'd42; b = 8'd170;  #10 
a = 8'd42; b = 8'd171;  #10 
a = 8'd42; b = 8'd172;  #10 
a = 8'd42; b = 8'd173;  #10 
a = 8'd42; b = 8'd174;  #10 
a = 8'd42; b = 8'd175;  #10 
a = 8'd42; b = 8'd176;  #10 
a = 8'd42; b = 8'd177;  #10 
a = 8'd42; b = 8'd178;  #10 
a = 8'd42; b = 8'd179;  #10 
a = 8'd42; b = 8'd180;  #10 
a = 8'd42; b = 8'd181;  #10 
a = 8'd42; b = 8'd182;  #10 
a = 8'd42; b = 8'd183;  #10 
a = 8'd42; b = 8'd184;  #10 
a = 8'd42; b = 8'd185;  #10 
a = 8'd42; b = 8'd186;  #10 
a = 8'd42; b = 8'd187;  #10 
a = 8'd42; b = 8'd188;  #10 
a = 8'd42; b = 8'd189;  #10 
a = 8'd42; b = 8'd190;  #10 
a = 8'd42; b = 8'd191;  #10 
a = 8'd42; b = 8'd192;  #10 
a = 8'd42; b = 8'd193;  #10 
a = 8'd42; b = 8'd194;  #10 
a = 8'd42; b = 8'd195;  #10 
a = 8'd42; b = 8'd196;  #10 
a = 8'd42; b = 8'd197;  #10 
a = 8'd42; b = 8'd198;  #10 
a = 8'd42; b = 8'd199;  #10 
a = 8'd42; b = 8'd200;  #10 
a = 8'd42; b = 8'd201;  #10 
a = 8'd42; b = 8'd202;  #10 
a = 8'd42; b = 8'd203;  #10 
a = 8'd42; b = 8'd204;  #10 
a = 8'd42; b = 8'd205;  #10 
a = 8'd42; b = 8'd206;  #10 
a = 8'd42; b = 8'd207;  #10 
a = 8'd42; b = 8'd208;  #10 
a = 8'd42; b = 8'd209;  #10 
a = 8'd42; b = 8'd210;  #10 
a = 8'd42; b = 8'd211;  #10 
a = 8'd42; b = 8'd212;  #10 
a = 8'd42; b = 8'd213;  #10 
a = 8'd42; b = 8'd214;  #10 
a = 8'd42; b = 8'd215;  #10 
a = 8'd42; b = 8'd216;  #10 
a = 8'd42; b = 8'd217;  #10 
a = 8'd42; b = 8'd218;  #10 
a = 8'd42; b = 8'd219;  #10 
a = 8'd42; b = 8'd220;  #10 
a = 8'd42; b = 8'd221;  #10 
a = 8'd42; b = 8'd222;  #10 
a = 8'd42; b = 8'd223;  #10 
a = 8'd42; b = 8'd224;  #10 
a = 8'd42; b = 8'd225;  #10 
a = 8'd42; b = 8'd226;  #10 
a = 8'd42; b = 8'd227;  #10 
a = 8'd42; b = 8'd228;  #10 
a = 8'd42; b = 8'd229;  #10 
a = 8'd42; b = 8'd230;  #10 
a = 8'd42; b = 8'd231;  #10 
a = 8'd42; b = 8'd232;  #10 
a = 8'd42; b = 8'd233;  #10 
a = 8'd42; b = 8'd234;  #10 
a = 8'd42; b = 8'd235;  #10 
a = 8'd42; b = 8'd236;  #10 
a = 8'd42; b = 8'd237;  #10 
a = 8'd42; b = 8'd238;  #10 
a = 8'd42; b = 8'd239;  #10 
a = 8'd42; b = 8'd240;  #10 
a = 8'd42; b = 8'd241;  #10 
a = 8'd42; b = 8'd242;  #10 
a = 8'd42; b = 8'd243;  #10 
a = 8'd42; b = 8'd244;  #10 
a = 8'd42; b = 8'd245;  #10 
a = 8'd42; b = 8'd246;  #10 
a = 8'd42; b = 8'd247;  #10 
a = 8'd42; b = 8'd248;  #10 
a = 8'd42; b = 8'd249;  #10 
a = 8'd42; b = 8'd250;  #10 
a = 8'd42; b = 8'd251;  #10 
a = 8'd42; b = 8'd252;  #10 
a = 8'd42; b = 8'd253;  #10 
a = 8'd42; b = 8'd254;  #10 
a = 8'd42; b = 8'd255;  #10 
a = 8'd43; b = 8'd0;  #10 
a = 8'd43; b = 8'd1;  #10 
a = 8'd43; b = 8'd2;  #10 
a = 8'd43; b = 8'd3;  #10 
a = 8'd43; b = 8'd4;  #10 
a = 8'd43; b = 8'd5;  #10 
a = 8'd43; b = 8'd6;  #10 
a = 8'd43; b = 8'd7;  #10 
a = 8'd43; b = 8'd8;  #10 
a = 8'd43; b = 8'd9;  #10 
a = 8'd43; b = 8'd10;  #10 
a = 8'd43; b = 8'd11;  #10 
a = 8'd43; b = 8'd12;  #10 
a = 8'd43; b = 8'd13;  #10 
a = 8'd43; b = 8'd14;  #10 
a = 8'd43; b = 8'd15;  #10 
a = 8'd43; b = 8'd16;  #10 
a = 8'd43; b = 8'd17;  #10 
a = 8'd43; b = 8'd18;  #10 
a = 8'd43; b = 8'd19;  #10 
a = 8'd43; b = 8'd20;  #10 
a = 8'd43; b = 8'd21;  #10 
a = 8'd43; b = 8'd22;  #10 
a = 8'd43; b = 8'd23;  #10 
a = 8'd43; b = 8'd24;  #10 
a = 8'd43; b = 8'd25;  #10 
a = 8'd43; b = 8'd26;  #10 
a = 8'd43; b = 8'd27;  #10 
a = 8'd43; b = 8'd28;  #10 
a = 8'd43; b = 8'd29;  #10 
a = 8'd43; b = 8'd30;  #10 
a = 8'd43; b = 8'd31;  #10 
a = 8'd43; b = 8'd32;  #10 
a = 8'd43; b = 8'd33;  #10 
a = 8'd43; b = 8'd34;  #10 
a = 8'd43; b = 8'd35;  #10 
a = 8'd43; b = 8'd36;  #10 
a = 8'd43; b = 8'd37;  #10 
a = 8'd43; b = 8'd38;  #10 
a = 8'd43; b = 8'd39;  #10 
a = 8'd43; b = 8'd40;  #10 
a = 8'd43; b = 8'd41;  #10 
a = 8'd43; b = 8'd42;  #10 
a = 8'd43; b = 8'd43;  #10 
a = 8'd43; b = 8'd44;  #10 
a = 8'd43; b = 8'd45;  #10 
a = 8'd43; b = 8'd46;  #10 
a = 8'd43; b = 8'd47;  #10 
a = 8'd43; b = 8'd48;  #10 
a = 8'd43; b = 8'd49;  #10 
a = 8'd43; b = 8'd50;  #10 
a = 8'd43; b = 8'd51;  #10 
a = 8'd43; b = 8'd52;  #10 
a = 8'd43; b = 8'd53;  #10 
a = 8'd43; b = 8'd54;  #10 
a = 8'd43; b = 8'd55;  #10 
a = 8'd43; b = 8'd56;  #10 
a = 8'd43; b = 8'd57;  #10 
a = 8'd43; b = 8'd58;  #10 
a = 8'd43; b = 8'd59;  #10 
a = 8'd43; b = 8'd60;  #10 
a = 8'd43; b = 8'd61;  #10 
a = 8'd43; b = 8'd62;  #10 
a = 8'd43; b = 8'd63;  #10 
a = 8'd43; b = 8'd64;  #10 
a = 8'd43; b = 8'd65;  #10 
a = 8'd43; b = 8'd66;  #10 
a = 8'd43; b = 8'd67;  #10 
a = 8'd43; b = 8'd68;  #10 
a = 8'd43; b = 8'd69;  #10 
a = 8'd43; b = 8'd70;  #10 
a = 8'd43; b = 8'd71;  #10 
a = 8'd43; b = 8'd72;  #10 
a = 8'd43; b = 8'd73;  #10 
a = 8'd43; b = 8'd74;  #10 
a = 8'd43; b = 8'd75;  #10 
a = 8'd43; b = 8'd76;  #10 
a = 8'd43; b = 8'd77;  #10 
a = 8'd43; b = 8'd78;  #10 
a = 8'd43; b = 8'd79;  #10 
a = 8'd43; b = 8'd80;  #10 
a = 8'd43; b = 8'd81;  #10 
a = 8'd43; b = 8'd82;  #10 
a = 8'd43; b = 8'd83;  #10 
a = 8'd43; b = 8'd84;  #10 
a = 8'd43; b = 8'd85;  #10 
a = 8'd43; b = 8'd86;  #10 
a = 8'd43; b = 8'd87;  #10 
a = 8'd43; b = 8'd88;  #10 
a = 8'd43; b = 8'd89;  #10 
a = 8'd43; b = 8'd90;  #10 
a = 8'd43; b = 8'd91;  #10 
a = 8'd43; b = 8'd92;  #10 
a = 8'd43; b = 8'd93;  #10 
a = 8'd43; b = 8'd94;  #10 
a = 8'd43; b = 8'd95;  #10 
a = 8'd43; b = 8'd96;  #10 
a = 8'd43; b = 8'd97;  #10 
a = 8'd43; b = 8'd98;  #10 
a = 8'd43; b = 8'd99;  #10 
a = 8'd43; b = 8'd100;  #10 
a = 8'd43; b = 8'd101;  #10 
a = 8'd43; b = 8'd102;  #10 
a = 8'd43; b = 8'd103;  #10 
a = 8'd43; b = 8'd104;  #10 
a = 8'd43; b = 8'd105;  #10 
a = 8'd43; b = 8'd106;  #10 
a = 8'd43; b = 8'd107;  #10 
a = 8'd43; b = 8'd108;  #10 
a = 8'd43; b = 8'd109;  #10 
a = 8'd43; b = 8'd110;  #10 
a = 8'd43; b = 8'd111;  #10 
a = 8'd43; b = 8'd112;  #10 
a = 8'd43; b = 8'd113;  #10 
a = 8'd43; b = 8'd114;  #10 
a = 8'd43; b = 8'd115;  #10 
a = 8'd43; b = 8'd116;  #10 
a = 8'd43; b = 8'd117;  #10 
a = 8'd43; b = 8'd118;  #10 
a = 8'd43; b = 8'd119;  #10 
a = 8'd43; b = 8'd120;  #10 
a = 8'd43; b = 8'd121;  #10 
a = 8'd43; b = 8'd122;  #10 
a = 8'd43; b = 8'd123;  #10 
a = 8'd43; b = 8'd124;  #10 
a = 8'd43; b = 8'd125;  #10 
a = 8'd43; b = 8'd126;  #10 
a = 8'd43; b = 8'd127;  #10 
a = 8'd43; b = 8'd128;  #10 
a = 8'd43; b = 8'd129;  #10 
a = 8'd43; b = 8'd130;  #10 
a = 8'd43; b = 8'd131;  #10 
a = 8'd43; b = 8'd132;  #10 
a = 8'd43; b = 8'd133;  #10 
a = 8'd43; b = 8'd134;  #10 
a = 8'd43; b = 8'd135;  #10 
a = 8'd43; b = 8'd136;  #10 
a = 8'd43; b = 8'd137;  #10 
a = 8'd43; b = 8'd138;  #10 
a = 8'd43; b = 8'd139;  #10 
a = 8'd43; b = 8'd140;  #10 
a = 8'd43; b = 8'd141;  #10 
a = 8'd43; b = 8'd142;  #10 
a = 8'd43; b = 8'd143;  #10 
a = 8'd43; b = 8'd144;  #10 
a = 8'd43; b = 8'd145;  #10 
a = 8'd43; b = 8'd146;  #10 
a = 8'd43; b = 8'd147;  #10 
a = 8'd43; b = 8'd148;  #10 
a = 8'd43; b = 8'd149;  #10 
a = 8'd43; b = 8'd150;  #10 
a = 8'd43; b = 8'd151;  #10 
a = 8'd43; b = 8'd152;  #10 
a = 8'd43; b = 8'd153;  #10 
a = 8'd43; b = 8'd154;  #10 
a = 8'd43; b = 8'd155;  #10 
a = 8'd43; b = 8'd156;  #10 
a = 8'd43; b = 8'd157;  #10 
a = 8'd43; b = 8'd158;  #10 
a = 8'd43; b = 8'd159;  #10 
a = 8'd43; b = 8'd160;  #10 
a = 8'd43; b = 8'd161;  #10 
a = 8'd43; b = 8'd162;  #10 
a = 8'd43; b = 8'd163;  #10 
a = 8'd43; b = 8'd164;  #10 
a = 8'd43; b = 8'd165;  #10 
a = 8'd43; b = 8'd166;  #10 
a = 8'd43; b = 8'd167;  #10 
a = 8'd43; b = 8'd168;  #10 
a = 8'd43; b = 8'd169;  #10 
a = 8'd43; b = 8'd170;  #10 
a = 8'd43; b = 8'd171;  #10 
a = 8'd43; b = 8'd172;  #10 
a = 8'd43; b = 8'd173;  #10 
a = 8'd43; b = 8'd174;  #10 
a = 8'd43; b = 8'd175;  #10 
a = 8'd43; b = 8'd176;  #10 
a = 8'd43; b = 8'd177;  #10 
a = 8'd43; b = 8'd178;  #10 
a = 8'd43; b = 8'd179;  #10 
a = 8'd43; b = 8'd180;  #10 
a = 8'd43; b = 8'd181;  #10 
a = 8'd43; b = 8'd182;  #10 
a = 8'd43; b = 8'd183;  #10 
a = 8'd43; b = 8'd184;  #10 
a = 8'd43; b = 8'd185;  #10 
a = 8'd43; b = 8'd186;  #10 
a = 8'd43; b = 8'd187;  #10 
a = 8'd43; b = 8'd188;  #10 
a = 8'd43; b = 8'd189;  #10 
a = 8'd43; b = 8'd190;  #10 
a = 8'd43; b = 8'd191;  #10 
a = 8'd43; b = 8'd192;  #10 
a = 8'd43; b = 8'd193;  #10 
a = 8'd43; b = 8'd194;  #10 
a = 8'd43; b = 8'd195;  #10 
a = 8'd43; b = 8'd196;  #10 
a = 8'd43; b = 8'd197;  #10 
a = 8'd43; b = 8'd198;  #10 
a = 8'd43; b = 8'd199;  #10 
a = 8'd43; b = 8'd200;  #10 
a = 8'd43; b = 8'd201;  #10 
a = 8'd43; b = 8'd202;  #10 
a = 8'd43; b = 8'd203;  #10 
a = 8'd43; b = 8'd204;  #10 
a = 8'd43; b = 8'd205;  #10 
a = 8'd43; b = 8'd206;  #10 
a = 8'd43; b = 8'd207;  #10 
a = 8'd43; b = 8'd208;  #10 
a = 8'd43; b = 8'd209;  #10 
a = 8'd43; b = 8'd210;  #10 
a = 8'd43; b = 8'd211;  #10 
a = 8'd43; b = 8'd212;  #10 
a = 8'd43; b = 8'd213;  #10 
a = 8'd43; b = 8'd214;  #10 
a = 8'd43; b = 8'd215;  #10 
a = 8'd43; b = 8'd216;  #10 
a = 8'd43; b = 8'd217;  #10 
a = 8'd43; b = 8'd218;  #10 
a = 8'd43; b = 8'd219;  #10 
a = 8'd43; b = 8'd220;  #10 
a = 8'd43; b = 8'd221;  #10 
a = 8'd43; b = 8'd222;  #10 
a = 8'd43; b = 8'd223;  #10 
a = 8'd43; b = 8'd224;  #10 
a = 8'd43; b = 8'd225;  #10 
a = 8'd43; b = 8'd226;  #10 
a = 8'd43; b = 8'd227;  #10 
a = 8'd43; b = 8'd228;  #10 
a = 8'd43; b = 8'd229;  #10 
a = 8'd43; b = 8'd230;  #10 
a = 8'd43; b = 8'd231;  #10 
a = 8'd43; b = 8'd232;  #10 
a = 8'd43; b = 8'd233;  #10 
a = 8'd43; b = 8'd234;  #10 
a = 8'd43; b = 8'd235;  #10 
a = 8'd43; b = 8'd236;  #10 
a = 8'd43; b = 8'd237;  #10 
a = 8'd43; b = 8'd238;  #10 
a = 8'd43; b = 8'd239;  #10 
a = 8'd43; b = 8'd240;  #10 
a = 8'd43; b = 8'd241;  #10 
a = 8'd43; b = 8'd242;  #10 
a = 8'd43; b = 8'd243;  #10 
a = 8'd43; b = 8'd244;  #10 
a = 8'd43; b = 8'd245;  #10 
a = 8'd43; b = 8'd246;  #10 
a = 8'd43; b = 8'd247;  #10 
a = 8'd43; b = 8'd248;  #10 
a = 8'd43; b = 8'd249;  #10 
a = 8'd43; b = 8'd250;  #10 
a = 8'd43; b = 8'd251;  #10 
a = 8'd43; b = 8'd252;  #10 
a = 8'd43; b = 8'd253;  #10 
a = 8'd43; b = 8'd254;  #10 
a = 8'd43; b = 8'd255;  #10 
a = 8'd44; b = 8'd0;  #10 
a = 8'd44; b = 8'd1;  #10 
a = 8'd44; b = 8'd2;  #10 
a = 8'd44; b = 8'd3;  #10 
a = 8'd44; b = 8'd4;  #10 
a = 8'd44; b = 8'd5;  #10 
a = 8'd44; b = 8'd6;  #10 
a = 8'd44; b = 8'd7;  #10 
a = 8'd44; b = 8'd8;  #10 
a = 8'd44; b = 8'd9;  #10 
a = 8'd44; b = 8'd10;  #10 
a = 8'd44; b = 8'd11;  #10 
a = 8'd44; b = 8'd12;  #10 
a = 8'd44; b = 8'd13;  #10 
a = 8'd44; b = 8'd14;  #10 
a = 8'd44; b = 8'd15;  #10 
a = 8'd44; b = 8'd16;  #10 
a = 8'd44; b = 8'd17;  #10 
a = 8'd44; b = 8'd18;  #10 
a = 8'd44; b = 8'd19;  #10 
a = 8'd44; b = 8'd20;  #10 
a = 8'd44; b = 8'd21;  #10 
a = 8'd44; b = 8'd22;  #10 
a = 8'd44; b = 8'd23;  #10 
a = 8'd44; b = 8'd24;  #10 
a = 8'd44; b = 8'd25;  #10 
a = 8'd44; b = 8'd26;  #10 
a = 8'd44; b = 8'd27;  #10 
a = 8'd44; b = 8'd28;  #10 
a = 8'd44; b = 8'd29;  #10 
a = 8'd44; b = 8'd30;  #10 
a = 8'd44; b = 8'd31;  #10 
a = 8'd44; b = 8'd32;  #10 
a = 8'd44; b = 8'd33;  #10 
a = 8'd44; b = 8'd34;  #10 
a = 8'd44; b = 8'd35;  #10 
a = 8'd44; b = 8'd36;  #10 
a = 8'd44; b = 8'd37;  #10 
a = 8'd44; b = 8'd38;  #10 
a = 8'd44; b = 8'd39;  #10 
a = 8'd44; b = 8'd40;  #10 
a = 8'd44; b = 8'd41;  #10 
a = 8'd44; b = 8'd42;  #10 
a = 8'd44; b = 8'd43;  #10 
a = 8'd44; b = 8'd44;  #10 
a = 8'd44; b = 8'd45;  #10 
a = 8'd44; b = 8'd46;  #10 
a = 8'd44; b = 8'd47;  #10 
a = 8'd44; b = 8'd48;  #10 
a = 8'd44; b = 8'd49;  #10 
a = 8'd44; b = 8'd50;  #10 
a = 8'd44; b = 8'd51;  #10 
a = 8'd44; b = 8'd52;  #10 
a = 8'd44; b = 8'd53;  #10 
a = 8'd44; b = 8'd54;  #10 
a = 8'd44; b = 8'd55;  #10 
a = 8'd44; b = 8'd56;  #10 
a = 8'd44; b = 8'd57;  #10 
a = 8'd44; b = 8'd58;  #10 
a = 8'd44; b = 8'd59;  #10 
a = 8'd44; b = 8'd60;  #10 
a = 8'd44; b = 8'd61;  #10 
a = 8'd44; b = 8'd62;  #10 
a = 8'd44; b = 8'd63;  #10 
a = 8'd44; b = 8'd64;  #10 
a = 8'd44; b = 8'd65;  #10 
a = 8'd44; b = 8'd66;  #10 
a = 8'd44; b = 8'd67;  #10 
a = 8'd44; b = 8'd68;  #10 
a = 8'd44; b = 8'd69;  #10 
a = 8'd44; b = 8'd70;  #10 
a = 8'd44; b = 8'd71;  #10 
a = 8'd44; b = 8'd72;  #10 
a = 8'd44; b = 8'd73;  #10 
a = 8'd44; b = 8'd74;  #10 
a = 8'd44; b = 8'd75;  #10 
a = 8'd44; b = 8'd76;  #10 
a = 8'd44; b = 8'd77;  #10 
a = 8'd44; b = 8'd78;  #10 
a = 8'd44; b = 8'd79;  #10 
a = 8'd44; b = 8'd80;  #10 
a = 8'd44; b = 8'd81;  #10 
a = 8'd44; b = 8'd82;  #10 
a = 8'd44; b = 8'd83;  #10 
a = 8'd44; b = 8'd84;  #10 
a = 8'd44; b = 8'd85;  #10 
a = 8'd44; b = 8'd86;  #10 
a = 8'd44; b = 8'd87;  #10 
a = 8'd44; b = 8'd88;  #10 
a = 8'd44; b = 8'd89;  #10 
a = 8'd44; b = 8'd90;  #10 
a = 8'd44; b = 8'd91;  #10 
a = 8'd44; b = 8'd92;  #10 
a = 8'd44; b = 8'd93;  #10 
a = 8'd44; b = 8'd94;  #10 
a = 8'd44; b = 8'd95;  #10 
a = 8'd44; b = 8'd96;  #10 
a = 8'd44; b = 8'd97;  #10 
a = 8'd44; b = 8'd98;  #10 
a = 8'd44; b = 8'd99;  #10 
a = 8'd44; b = 8'd100;  #10 
a = 8'd44; b = 8'd101;  #10 
a = 8'd44; b = 8'd102;  #10 
a = 8'd44; b = 8'd103;  #10 
a = 8'd44; b = 8'd104;  #10 
a = 8'd44; b = 8'd105;  #10 
a = 8'd44; b = 8'd106;  #10 
a = 8'd44; b = 8'd107;  #10 
a = 8'd44; b = 8'd108;  #10 
a = 8'd44; b = 8'd109;  #10 
a = 8'd44; b = 8'd110;  #10 
a = 8'd44; b = 8'd111;  #10 
a = 8'd44; b = 8'd112;  #10 
a = 8'd44; b = 8'd113;  #10 
a = 8'd44; b = 8'd114;  #10 
a = 8'd44; b = 8'd115;  #10 
a = 8'd44; b = 8'd116;  #10 
a = 8'd44; b = 8'd117;  #10 
a = 8'd44; b = 8'd118;  #10 
a = 8'd44; b = 8'd119;  #10 
a = 8'd44; b = 8'd120;  #10 
a = 8'd44; b = 8'd121;  #10 
a = 8'd44; b = 8'd122;  #10 
a = 8'd44; b = 8'd123;  #10 
a = 8'd44; b = 8'd124;  #10 
a = 8'd44; b = 8'd125;  #10 
a = 8'd44; b = 8'd126;  #10 
a = 8'd44; b = 8'd127;  #10 
a = 8'd44; b = 8'd128;  #10 
a = 8'd44; b = 8'd129;  #10 
a = 8'd44; b = 8'd130;  #10 
a = 8'd44; b = 8'd131;  #10 
a = 8'd44; b = 8'd132;  #10 
a = 8'd44; b = 8'd133;  #10 
a = 8'd44; b = 8'd134;  #10 
a = 8'd44; b = 8'd135;  #10 
a = 8'd44; b = 8'd136;  #10 
a = 8'd44; b = 8'd137;  #10 
a = 8'd44; b = 8'd138;  #10 
a = 8'd44; b = 8'd139;  #10 
a = 8'd44; b = 8'd140;  #10 
a = 8'd44; b = 8'd141;  #10 
a = 8'd44; b = 8'd142;  #10 
a = 8'd44; b = 8'd143;  #10 
a = 8'd44; b = 8'd144;  #10 
a = 8'd44; b = 8'd145;  #10 
a = 8'd44; b = 8'd146;  #10 
a = 8'd44; b = 8'd147;  #10 
a = 8'd44; b = 8'd148;  #10 
a = 8'd44; b = 8'd149;  #10 
a = 8'd44; b = 8'd150;  #10 
a = 8'd44; b = 8'd151;  #10 
a = 8'd44; b = 8'd152;  #10 
a = 8'd44; b = 8'd153;  #10 
a = 8'd44; b = 8'd154;  #10 
a = 8'd44; b = 8'd155;  #10 
a = 8'd44; b = 8'd156;  #10 
a = 8'd44; b = 8'd157;  #10 
a = 8'd44; b = 8'd158;  #10 
a = 8'd44; b = 8'd159;  #10 
a = 8'd44; b = 8'd160;  #10 
a = 8'd44; b = 8'd161;  #10 
a = 8'd44; b = 8'd162;  #10 
a = 8'd44; b = 8'd163;  #10 
a = 8'd44; b = 8'd164;  #10 
a = 8'd44; b = 8'd165;  #10 
a = 8'd44; b = 8'd166;  #10 
a = 8'd44; b = 8'd167;  #10 
a = 8'd44; b = 8'd168;  #10 
a = 8'd44; b = 8'd169;  #10 
a = 8'd44; b = 8'd170;  #10 
a = 8'd44; b = 8'd171;  #10 
a = 8'd44; b = 8'd172;  #10 
a = 8'd44; b = 8'd173;  #10 
a = 8'd44; b = 8'd174;  #10 
a = 8'd44; b = 8'd175;  #10 
a = 8'd44; b = 8'd176;  #10 
a = 8'd44; b = 8'd177;  #10 
a = 8'd44; b = 8'd178;  #10 
a = 8'd44; b = 8'd179;  #10 
a = 8'd44; b = 8'd180;  #10 
a = 8'd44; b = 8'd181;  #10 
a = 8'd44; b = 8'd182;  #10 
a = 8'd44; b = 8'd183;  #10 
a = 8'd44; b = 8'd184;  #10 
a = 8'd44; b = 8'd185;  #10 
a = 8'd44; b = 8'd186;  #10 
a = 8'd44; b = 8'd187;  #10 
a = 8'd44; b = 8'd188;  #10 
a = 8'd44; b = 8'd189;  #10 
a = 8'd44; b = 8'd190;  #10 
a = 8'd44; b = 8'd191;  #10 
a = 8'd44; b = 8'd192;  #10 
a = 8'd44; b = 8'd193;  #10 
a = 8'd44; b = 8'd194;  #10 
a = 8'd44; b = 8'd195;  #10 
a = 8'd44; b = 8'd196;  #10 
a = 8'd44; b = 8'd197;  #10 
a = 8'd44; b = 8'd198;  #10 
a = 8'd44; b = 8'd199;  #10 
a = 8'd44; b = 8'd200;  #10 
a = 8'd44; b = 8'd201;  #10 
a = 8'd44; b = 8'd202;  #10 
a = 8'd44; b = 8'd203;  #10 
a = 8'd44; b = 8'd204;  #10 
a = 8'd44; b = 8'd205;  #10 
a = 8'd44; b = 8'd206;  #10 
a = 8'd44; b = 8'd207;  #10 
a = 8'd44; b = 8'd208;  #10 
a = 8'd44; b = 8'd209;  #10 
a = 8'd44; b = 8'd210;  #10 
a = 8'd44; b = 8'd211;  #10 
a = 8'd44; b = 8'd212;  #10 
a = 8'd44; b = 8'd213;  #10 
a = 8'd44; b = 8'd214;  #10 
a = 8'd44; b = 8'd215;  #10 
a = 8'd44; b = 8'd216;  #10 
a = 8'd44; b = 8'd217;  #10 
a = 8'd44; b = 8'd218;  #10 
a = 8'd44; b = 8'd219;  #10 
a = 8'd44; b = 8'd220;  #10 
a = 8'd44; b = 8'd221;  #10 
a = 8'd44; b = 8'd222;  #10 
a = 8'd44; b = 8'd223;  #10 
a = 8'd44; b = 8'd224;  #10 
a = 8'd44; b = 8'd225;  #10 
a = 8'd44; b = 8'd226;  #10 
a = 8'd44; b = 8'd227;  #10 
a = 8'd44; b = 8'd228;  #10 
a = 8'd44; b = 8'd229;  #10 
a = 8'd44; b = 8'd230;  #10 
a = 8'd44; b = 8'd231;  #10 
a = 8'd44; b = 8'd232;  #10 
a = 8'd44; b = 8'd233;  #10 
a = 8'd44; b = 8'd234;  #10 
a = 8'd44; b = 8'd235;  #10 
a = 8'd44; b = 8'd236;  #10 
a = 8'd44; b = 8'd237;  #10 
a = 8'd44; b = 8'd238;  #10 
a = 8'd44; b = 8'd239;  #10 
a = 8'd44; b = 8'd240;  #10 
a = 8'd44; b = 8'd241;  #10 
a = 8'd44; b = 8'd242;  #10 
a = 8'd44; b = 8'd243;  #10 
a = 8'd44; b = 8'd244;  #10 
a = 8'd44; b = 8'd245;  #10 
a = 8'd44; b = 8'd246;  #10 
a = 8'd44; b = 8'd247;  #10 
a = 8'd44; b = 8'd248;  #10 
a = 8'd44; b = 8'd249;  #10 
a = 8'd44; b = 8'd250;  #10 
a = 8'd44; b = 8'd251;  #10 
a = 8'd44; b = 8'd252;  #10 
a = 8'd44; b = 8'd253;  #10 
a = 8'd44; b = 8'd254;  #10 
a = 8'd44; b = 8'd255;  #10 
a = 8'd45; b = 8'd0;  #10 
a = 8'd45; b = 8'd1;  #10 
a = 8'd45; b = 8'd2;  #10 
a = 8'd45; b = 8'd3;  #10 
a = 8'd45; b = 8'd4;  #10 
a = 8'd45; b = 8'd5;  #10 
a = 8'd45; b = 8'd6;  #10 
a = 8'd45; b = 8'd7;  #10 
a = 8'd45; b = 8'd8;  #10 
a = 8'd45; b = 8'd9;  #10 
a = 8'd45; b = 8'd10;  #10 
a = 8'd45; b = 8'd11;  #10 
a = 8'd45; b = 8'd12;  #10 
a = 8'd45; b = 8'd13;  #10 
a = 8'd45; b = 8'd14;  #10 
a = 8'd45; b = 8'd15;  #10 
a = 8'd45; b = 8'd16;  #10 
a = 8'd45; b = 8'd17;  #10 
a = 8'd45; b = 8'd18;  #10 
a = 8'd45; b = 8'd19;  #10 
a = 8'd45; b = 8'd20;  #10 
a = 8'd45; b = 8'd21;  #10 
a = 8'd45; b = 8'd22;  #10 
a = 8'd45; b = 8'd23;  #10 
a = 8'd45; b = 8'd24;  #10 
a = 8'd45; b = 8'd25;  #10 
a = 8'd45; b = 8'd26;  #10 
a = 8'd45; b = 8'd27;  #10 
a = 8'd45; b = 8'd28;  #10 
a = 8'd45; b = 8'd29;  #10 
a = 8'd45; b = 8'd30;  #10 
a = 8'd45; b = 8'd31;  #10 
a = 8'd45; b = 8'd32;  #10 
a = 8'd45; b = 8'd33;  #10 
a = 8'd45; b = 8'd34;  #10 
a = 8'd45; b = 8'd35;  #10 
a = 8'd45; b = 8'd36;  #10 
a = 8'd45; b = 8'd37;  #10 
a = 8'd45; b = 8'd38;  #10 
a = 8'd45; b = 8'd39;  #10 
a = 8'd45; b = 8'd40;  #10 
a = 8'd45; b = 8'd41;  #10 
a = 8'd45; b = 8'd42;  #10 
a = 8'd45; b = 8'd43;  #10 
a = 8'd45; b = 8'd44;  #10 
a = 8'd45; b = 8'd45;  #10 
a = 8'd45; b = 8'd46;  #10 
a = 8'd45; b = 8'd47;  #10 
a = 8'd45; b = 8'd48;  #10 
a = 8'd45; b = 8'd49;  #10 
a = 8'd45; b = 8'd50;  #10 
a = 8'd45; b = 8'd51;  #10 
a = 8'd45; b = 8'd52;  #10 
a = 8'd45; b = 8'd53;  #10 
a = 8'd45; b = 8'd54;  #10 
a = 8'd45; b = 8'd55;  #10 
a = 8'd45; b = 8'd56;  #10 
a = 8'd45; b = 8'd57;  #10 
a = 8'd45; b = 8'd58;  #10 
a = 8'd45; b = 8'd59;  #10 
a = 8'd45; b = 8'd60;  #10 
a = 8'd45; b = 8'd61;  #10 
a = 8'd45; b = 8'd62;  #10 
a = 8'd45; b = 8'd63;  #10 
a = 8'd45; b = 8'd64;  #10 
a = 8'd45; b = 8'd65;  #10 
a = 8'd45; b = 8'd66;  #10 
a = 8'd45; b = 8'd67;  #10 
a = 8'd45; b = 8'd68;  #10 
a = 8'd45; b = 8'd69;  #10 
a = 8'd45; b = 8'd70;  #10 
a = 8'd45; b = 8'd71;  #10 
a = 8'd45; b = 8'd72;  #10 
a = 8'd45; b = 8'd73;  #10 
a = 8'd45; b = 8'd74;  #10 
a = 8'd45; b = 8'd75;  #10 
a = 8'd45; b = 8'd76;  #10 
a = 8'd45; b = 8'd77;  #10 
a = 8'd45; b = 8'd78;  #10 
a = 8'd45; b = 8'd79;  #10 
a = 8'd45; b = 8'd80;  #10 
a = 8'd45; b = 8'd81;  #10 
a = 8'd45; b = 8'd82;  #10 
a = 8'd45; b = 8'd83;  #10 
a = 8'd45; b = 8'd84;  #10 
a = 8'd45; b = 8'd85;  #10 
a = 8'd45; b = 8'd86;  #10 
a = 8'd45; b = 8'd87;  #10 
a = 8'd45; b = 8'd88;  #10 
a = 8'd45; b = 8'd89;  #10 
a = 8'd45; b = 8'd90;  #10 
a = 8'd45; b = 8'd91;  #10 
a = 8'd45; b = 8'd92;  #10 
a = 8'd45; b = 8'd93;  #10 
a = 8'd45; b = 8'd94;  #10 
a = 8'd45; b = 8'd95;  #10 
a = 8'd45; b = 8'd96;  #10 
a = 8'd45; b = 8'd97;  #10 
a = 8'd45; b = 8'd98;  #10 
a = 8'd45; b = 8'd99;  #10 
a = 8'd45; b = 8'd100;  #10 
a = 8'd45; b = 8'd101;  #10 
a = 8'd45; b = 8'd102;  #10 
a = 8'd45; b = 8'd103;  #10 
a = 8'd45; b = 8'd104;  #10 
a = 8'd45; b = 8'd105;  #10 
a = 8'd45; b = 8'd106;  #10 
a = 8'd45; b = 8'd107;  #10 
a = 8'd45; b = 8'd108;  #10 
a = 8'd45; b = 8'd109;  #10 
a = 8'd45; b = 8'd110;  #10 
a = 8'd45; b = 8'd111;  #10 
a = 8'd45; b = 8'd112;  #10 
a = 8'd45; b = 8'd113;  #10 
a = 8'd45; b = 8'd114;  #10 
a = 8'd45; b = 8'd115;  #10 
a = 8'd45; b = 8'd116;  #10 
a = 8'd45; b = 8'd117;  #10 
a = 8'd45; b = 8'd118;  #10 
a = 8'd45; b = 8'd119;  #10 
a = 8'd45; b = 8'd120;  #10 
a = 8'd45; b = 8'd121;  #10 
a = 8'd45; b = 8'd122;  #10 
a = 8'd45; b = 8'd123;  #10 
a = 8'd45; b = 8'd124;  #10 
a = 8'd45; b = 8'd125;  #10 
a = 8'd45; b = 8'd126;  #10 
a = 8'd45; b = 8'd127;  #10 
a = 8'd45; b = 8'd128;  #10 
a = 8'd45; b = 8'd129;  #10 
a = 8'd45; b = 8'd130;  #10 
a = 8'd45; b = 8'd131;  #10 
a = 8'd45; b = 8'd132;  #10 
a = 8'd45; b = 8'd133;  #10 
a = 8'd45; b = 8'd134;  #10 
a = 8'd45; b = 8'd135;  #10 
a = 8'd45; b = 8'd136;  #10 
a = 8'd45; b = 8'd137;  #10 
a = 8'd45; b = 8'd138;  #10 
a = 8'd45; b = 8'd139;  #10 
a = 8'd45; b = 8'd140;  #10 
a = 8'd45; b = 8'd141;  #10 
a = 8'd45; b = 8'd142;  #10 
a = 8'd45; b = 8'd143;  #10 
a = 8'd45; b = 8'd144;  #10 
a = 8'd45; b = 8'd145;  #10 
a = 8'd45; b = 8'd146;  #10 
a = 8'd45; b = 8'd147;  #10 
a = 8'd45; b = 8'd148;  #10 
a = 8'd45; b = 8'd149;  #10 
a = 8'd45; b = 8'd150;  #10 
a = 8'd45; b = 8'd151;  #10 
a = 8'd45; b = 8'd152;  #10 
a = 8'd45; b = 8'd153;  #10 
a = 8'd45; b = 8'd154;  #10 
a = 8'd45; b = 8'd155;  #10 
a = 8'd45; b = 8'd156;  #10 
a = 8'd45; b = 8'd157;  #10 
a = 8'd45; b = 8'd158;  #10 
a = 8'd45; b = 8'd159;  #10 
a = 8'd45; b = 8'd160;  #10 
a = 8'd45; b = 8'd161;  #10 
a = 8'd45; b = 8'd162;  #10 
a = 8'd45; b = 8'd163;  #10 
a = 8'd45; b = 8'd164;  #10 
a = 8'd45; b = 8'd165;  #10 
a = 8'd45; b = 8'd166;  #10 
a = 8'd45; b = 8'd167;  #10 
a = 8'd45; b = 8'd168;  #10 
a = 8'd45; b = 8'd169;  #10 
a = 8'd45; b = 8'd170;  #10 
a = 8'd45; b = 8'd171;  #10 
a = 8'd45; b = 8'd172;  #10 
a = 8'd45; b = 8'd173;  #10 
a = 8'd45; b = 8'd174;  #10 
a = 8'd45; b = 8'd175;  #10 
a = 8'd45; b = 8'd176;  #10 
a = 8'd45; b = 8'd177;  #10 
a = 8'd45; b = 8'd178;  #10 
a = 8'd45; b = 8'd179;  #10 
a = 8'd45; b = 8'd180;  #10 
a = 8'd45; b = 8'd181;  #10 
a = 8'd45; b = 8'd182;  #10 
a = 8'd45; b = 8'd183;  #10 
a = 8'd45; b = 8'd184;  #10 
a = 8'd45; b = 8'd185;  #10 
a = 8'd45; b = 8'd186;  #10 
a = 8'd45; b = 8'd187;  #10 
a = 8'd45; b = 8'd188;  #10 
a = 8'd45; b = 8'd189;  #10 
a = 8'd45; b = 8'd190;  #10 
a = 8'd45; b = 8'd191;  #10 
a = 8'd45; b = 8'd192;  #10 
a = 8'd45; b = 8'd193;  #10 
a = 8'd45; b = 8'd194;  #10 
a = 8'd45; b = 8'd195;  #10 
a = 8'd45; b = 8'd196;  #10 
a = 8'd45; b = 8'd197;  #10 
a = 8'd45; b = 8'd198;  #10 
a = 8'd45; b = 8'd199;  #10 
a = 8'd45; b = 8'd200;  #10 
a = 8'd45; b = 8'd201;  #10 
a = 8'd45; b = 8'd202;  #10 
a = 8'd45; b = 8'd203;  #10 
a = 8'd45; b = 8'd204;  #10 
a = 8'd45; b = 8'd205;  #10 
a = 8'd45; b = 8'd206;  #10 
a = 8'd45; b = 8'd207;  #10 
a = 8'd45; b = 8'd208;  #10 
a = 8'd45; b = 8'd209;  #10 
a = 8'd45; b = 8'd210;  #10 
a = 8'd45; b = 8'd211;  #10 
a = 8'd45; b = 8'd212;  #10 
a = 8'd45; b = 8'd213;  #10 
a = 8'd45; b = 8'd214;  #10 
a = 8'd45; b = 8'd215;  #10 
a = 8'd45; b = 8'd216;  #10 
a = 8'd45; b = 8'd217;  #10 
a = 8'd45; b = 8'd218;  #10 
a = 8'd45; b = 8'd219;  #10 
a = 8'd45; b = 8'd220;  #10 
a = 8'd45; b = 8'd221;  #10 
a = 8'd45; b = 8'd222;  #10 
a = 8'd45; b = 8'd223;  #10 
a = 8'd45; b = 8'd224;  #10 
a = 8'd45; b = 8'd225;  #10 
a = 8'd45; b = 8'd226;  #10 
a = 8'd45; b = 8'd227;  #10 
a = 8'd45; b = 8'd228;  #10 
a = 8'd45; b = 8'd229;  #10 
a = 8'd45; b = 8'd230;  #10 
a = 8'd45; b = 8'd231;  #10 
a = 8'd45; b = 8'd232;  #10 
a = 8'd45; b = 8'd233;  #10 
a = 8'd45; b = 8'd234;  #10 
a = 8'd45; b = 8'd235;  #10 
a = 8'd45; b = 8'd236;  #10 
a = 8'd45; b = 8'd237;  #10 
a = 8'd45; b = 8'd238;  #10 
a = 8'd45; b = 8'd239;  #10 
a = 8'd45; b = 8'd240;  #10 
a = 8'd45; b = 8'd241;  #10 
a = 8'd45; b = 8'd242;  #10 
a = 8'd45; b = 8'd243;  #10 
a = 8'd45; b = 8'd244;  #10 
a = 8'd45; b = 8'd245;  #10 
a = 8'd45; b = 8'd246;  #10 
a = 8'd45; b = 8'd247;  #10 
a = 8'd45; b = 8'd248;  #10 
a = 8'd45; b = 8'd249;  #10 
a = 8'd45; b = 8'd250;  #10 
a = 8'd45; b = 8'd251;  #10 
a = 8'd45; b = 8'd252;  #10 
a = 8'd45; b = 8'd253;  #10 
a = 8'd45; b = 8'd254;  #10 
a = 8'd45; b = 8'd255;  #10 
a = 8'd46; b = 8'd0;  #10 
a = 8'd46; b = 8'd1;  #10 
a = 8'd46; b = 8'd2;  #10 
a = 8'd46; b = 8'd3;  #10 
a = 8'd46; b = 8'd4;  #10 
a = 8'd46; b = 8'd5;  #10 
a = 8'd46; b = 8'd6;  #10 
a = 8'd46; b = 8'd7;  #10 
a = 8'd46; b = 8'd8;  #10 
a = 8'd46; b = 8'd9;  #10 
a = 8'd46; b = 8'd10;  #10 
a = 8'd46; b = 8'd11;  #10 
a = 8'd46; b = 8'd12;  #10 
a = 8'd46; b = 8'd13;  #10 
a = 8'd46; b = 8'd14;  #10 
a = 8'd46; b = 8'd15;  #10 
a = 8'd46; b = 8'd16;  #10 
a = 8'd46; b = 8'd17;  #10 
a = 8'd46; b = 8'd18;  #10 
a = 8'd46; b = 8'd19;  #10 
a = 8'd46; b = 8'd20;  #10 
a = 8'd46; b = 8'd21;  #10 
a = 8'd46; b = 8'd22;  #10 
a = 8'd46; b = 8'd23;  #10 
a = 8'd46; b = 8'd24;  #10 
a = 8'd46; b = 8'd25;  #10 
a = 8'd46; b = 8'd26;  #10 
a = 8'd46; b = 8'd27;  #10 
a = 8'd46; b = 8'd28;  #10 
a = 8'd46; b = 8'd29;  #10 
a = 8'd46; b = 8'd30;  #10 
a = 8'd46; b = 8'd31;  #10 
a = 8'd46; b = 8'd32;  #10 
a = 8'd46; b = 8'd33;  #10 
a = 8'd46; b = 8'd34;  #10 
a = 8'd46; b = 8'd35;  #10 
a = 8'd46; b = 8'd36;  #10 
a = 8'd46; b = 8'd37;  #10 
a = 8'd46; b = 8'd38;  #10 
a = 8'd46; b = 8'd39;  #10 
a = 8'd46; b = 8'd40;  #10 
a = 8'd46; b = 8'd41;  #10 
a = 8'd46; b = 8'd42;  #10 
a = 8'd46; b = 8'd43;  #10 
a = 8'd46; b = 8'd44;  #10 
a = 8'd46; b = 8'd45;  #10 
a = 8'd46; b = 8'd46;  #10 
a = 8'd46; b = 8'd47;  #10 
a = 8'd46; b = 8'd48;  #10 
a = 8'd46; b = 8'd49;  #10 
a = 8'd46; b = 8'd50;  #10 
a = 8'd46; b = 8'd51;  #10 
a = 8'd46; b = 8'd52;  #10 
a = 8'd46; b = 8'd53;  #10 
a = 8'd46; b = 8'd54;  #10 
a = 8'd46; b = 8'd55;  #10 
a = 8'd46; b = 8'd56;  #10 
a = 8'd46; b = 8'd57;  #10 
a = 8'd46; b = 8'd58;  #10 
a = 8'd46; b = 8'd59;  #10 
a = 8'd46; b = 8'd60;  #10 
a = 8'd46; b = 8'd61;  #10 
a = 8'd46; b = 8'd62;  #10 
a = 8'd46; b = 8'd63;  #10 
a = 8'd46; b = 8'd64;  #10 
a = 8'd46; b = 8'd65;  #10 
a = 8'd46; b = 8'd66;  #10 
a = 8'd46; b = 8'd67;  #10 
a = 8'd46; b = 8'd68;  #10 
a = 8'd46; b = 8'd69;  #10 
a = 8'd46; b = 8'd70;  #10 
a = 8'd46; b = 8'd71;  #10 
a = 8'd46; b = 8'd72;  #10 
a = 8'd46; b = 8'd73;  #10 
a = 8'd46; b = 8'd74;  #10 
a = 8'd46; b = 8'd75;  #10 
a = 8'd46; b = 8'd76;  #10 
a = 8'd46; b = 8'd77;  #10 
a = 8'd46; b = 8'd78;  #10 
a = 8'd46; b = 8'd79;  #10 
a = 8'd46; b = 8'd80;  #10 
a = 8'd46; b = 8'd81;  #10 
a = 8'd46; b = 8'd82;  #10 
a = 8'd46; b = 8'd83;  #10 
a = 8'd46; b = 8'd84;  #10 
a = 8'd46; b = 8'd85;  #10 
a = 8'd46; b = 8'd86;  #10 
a = 8'd46; b = 8'd87;  #10 
a = 8'd46; b = 8'd88;  #10 
a = 8'd46; b = 8'd89;  #10 
a = 8'd46; b = 8'd90;  #10 
a = 8'd46; b = 8'd91;  #10 
a = 8'd46; b = 8'd92;  #10 
a = 8'd46; b = 8'd93;  #10 
a = 8'd46; b = 8'd94;  #10 
a = 8'd46; b = 8'd95;  #10 
a = 8'd46; b = 8'd96;  #10 
a = 8'd46; b = 8'd97;  #10 
a = 8'd46; b = 8'd98;  #10 
a = 8'd46; b = 8'd99;  #10 
a = 8'd46; b = 8'd100;  #10 
a = 8'd46; b = 8'd101;  #10 
a = 8'd46; b = 8'd102;  #10 
a = 8'd46; b = 8'd103;  #10 
a = 8'd46; b = 8'd104;  #10 
a = 8'd46; b = 8'd105;  #10 
a = 8'd46; b = 8'd106;  #10 
a = 8'd46; b = 8'd107;  #10 
a = 8'd46; b = 8'd108;  #10 
a = 8'd46; b = 8'd109;  #10 
a = 8'd46; b = 8'd110;  #10 
a = 8'd46; b = 8'd111;  #10 
a = 8'd46; b = 8'd112;  #10 
a = 8'd46; b = 8'd113;  #10 
a = 8'd46; b = 8'd114;  #10 
a = 8'd46; b = 8'd115;  #10 
a = 8'd46; b = 8'd116;  #10 
a = 8'd46; b = 8'd117;  #10 
a = 8'd46; b = 8'd118;  #10 
a = 8'd46; b = 8'd119;  #10 
a = 8'd46; b = 8'd120;  #10 
a = 8'd46; b = 8'd121;  #10 
a = 8'd46; b = 8'd122;  #10 
a = 8'd46; b = 8'd123;  #10 
a = 8'd46; b = 8'd124;  #10 
a = 8'd46; b = 8'd125;  #10 
a = 8'd46; b = 8'd126;  #10 
a = 8'd46; b = 8'd127;  #10 
a = 8'd46; b = 8'd128;  #10 
a = 8'd46; b = 8'd129;  #10 
a = 8'd46; b = 8'd130;  #10 
a = 8'd46; b = 8'd131;  #10 
a = 8'd46; b = 8'd132;  #10 
a = 8'd46; b = 8'd133;  #10 
a = 8'd46; b = 8'd134;  #10 
a = 8'd46; b = 8'd135;  #10 
a = 8'd46; b = 8'd136;  #10 
a = 8'd46; b = 8'd137;  #10 
a = 8'd46; b = 8'd138;  #10 
a = 8'd46; b = 8'd139;  #10 
a = 8'd46; b = 8'd140;  #10 
a = 8'd46; b = 8'd141;  #10 
a = 8'd46; b = 8'd142;  #10 
a = 8'd46; b = 8'd143;  #10 
a = 8'd46; b = 8'd144;  #10 
a = 8'd46; b = 8'd145;  #10 
a = 8'd46; b = 8'd146;  #10 
a = 8'd46; b = 8'd147;  #10 
a = 8'd46; b = 8'd148;  #10 
a = 8'd46; b = 8'd149;  #10 
a = 8'd46; b = 8'd150;  #10 
a = 8'd46; b = 8'd151;  #10 
a = 8'd46; b = 8'd152;  #10 
a = 8'd46; b = 8'd153;  #10 
a = 8'd46; b = 8'd154;  #10 
a = 8'd46; b = 8'd155;  #10 
a = 8'd46; b = 8'd156;  #10 
a = 8'd46; b = 8'd157;  #10 
a = 8'd46; b = 8'd158;  #10 
a = 8'd46; b = 8'd159;  #10 
a = 8'd46; b = 8'd160;  #10 
a = 8'd46; b = 8'd161;  #10 
a = 8'd46; b = 8'd162;  #10 
a = 8'd46; b = 8'd163;  #10 
a = 8'd46; b = 8'd164;  #10 
a = 8'd46; b = 8'd165;  #10 
a = 8'd46; b = 8'd166;  #10 
a = 8'd46; b = 8'd167;  #10 
a = 8'd46; b = 8'd168;  #10 
a = 8'd46; b = 8'd169;  #10 
a = 8'd46; b = 8'd170;  #10 
a = 8'd46; b = 8'd171;  #10 
a = 8'd46; b = 8'd172;  #10 
a = 8'd46; b = 8'd173;  #10 
a = 8'd46; b = 8'd174;  #10 
a = 8'd46; b = 8'd175;  #10 
a = 8'd46; b = 8'd176;  #10 
a = 8'd46; b = 8'd177;  #10 
a = 8'd46; b = 8'd178;  #10 
a = 8'd46; b = 8'd179;  #10 
a = 8'd46; b = 8'd180;  #10 
a = 8'd46; b = 8'd181;  #10 
a = 8'd46; b = 8'd182;  #10 
a = 8'd46; b = 8'd183;  #10 
a = 8'd46; b = 8'd184;  #10 
a = 8'd46; b = 8'd185;  #10 
a = 8'd46; b = 8'd186;  #10 
a = 8'd46; b = 8'd187;  #10 
a = 8'd46; b = 8'd188;  #10 
a = 8'd46; b = 8'd189;  #10 
a = 8'd46; b = 8'd190;  #10 
a = 8'd46; b = 8'd191;  #10 
a = 8'd46; b = 8'd192;  #10 
a = 8'd46; b = 8'd193;  #10 
a = 8'd46; b = 8'd194;  #10 
a = 8'd46; b = 8'd195;  #10 
a = 8'd46; b = 8'd196;  #10 
a = 8'd46; b = 8'd197;  #10 
a = 8'd46; b = 8'd198;  #10 
a = 8'd46; b = 8'd199;  #10 
a = 8'd46; b = 8'd200;  #10 
a = 8'd46; b = 8'd201;  #10 
a = 8'd46; b = 8'd202;  #10 
a = 8'd46; b = 8'd203;  #10 
a = 8'd46; b = 8'd204;  #10 
a = 8'd46; b = 8'd205;  #10 
a = 8'd46; b = 8'd206;  #10 
a = 8'd46; b = 8'd207;  #10 
a = 8'd46; b = 8'd208;  #10 
a = 8'd46; b = 8'd209;  #10 
a = 8'd46; b = 8'd210;  #10 
a = 8'd46; b = 8'd211;  #10 
a = 8'd46; b = 8'd212;  #10 
a = 8'd46; b = 8'd213;  #10 
a = 8'd46; b = 8'd214;  #10 
a = 8'd46; b = 8'd215;  #10 
a = 8'd46; b = 8'd216;  #10 
a = 8'd46; b = 8'd217;  #10 
a = 8'd46; b = 8'd218;  #10 
a = 8'd46; b = 8'd219;  #10 
a = 8'd46; b = 8'd220;  #10 
a = 8'd46; b = 8'd221;  #10 
a = 8'd46; b = 8'd222;  #10 
a = 8'd46; b = 8'd223;  #10 
a = 8'd46; b = 8'd224;  #10 
a = 8'd46; b = 8'd225;  #10 
a = 8'd46; b = 8'd226;  #10 
a = 8'd46; b = 8'd227;  #10 
a = 8'd46; b = 8'd228;  #10 
a = 8'd46; b = 8'd229;  #10 
a = 8'd46; b = 8'd230;  #10 
a = 8'd46; b = 8'd231;  #10 
a = 8'd46; b = 8'd232;  #10 
a = 8'd46; b = 8'd233;  #10 
a = 8'd46; b = 8'd234;  #10 
a = 8'd46; b = 8'd235;  #10 
a = 8'd46; b = 8'd236;  #10 
a = 8'd46; b = 8'd237;  #10 
a = 8'd46; b = 8'd238;  #10 
a = 8'd46; b = 8'd239;  #10 
a = 8'd46; b = 8'd240;  #10 
a = 8'd46; b = 8'd241;  #10 
a = 8'd46; b = 8'd242;  #10 
a = 8'd46; b = 8'd243;  #10 
a = 8'd46; b = 8'd244;  #10 
a = 8'd46; b = 8'd245;  #10 
a = 8'd46; b = 8'd246;  #10 
a = 8'd46; b = 8'd247;  #10 
a = 8'd46; b = 8'd248;  #10 
a = 8'd46; b = 8'd249;  #10 
a = 8'd46; b = 8'd250;  #10 
a = 8'd46; b = 8'd251;  #10 
a = 8'd46; b = 8'd252;  #10 
a = 8'd46; b = 8'd253;  #10 
a = 8'd46; b = 8'd254;  #10 
a = 8'd46; b = 8'd255;  #10 
a = 8'd47; b = 8'd0;  #10 
a = 8'd47; b = 8'd1;  #10 
a = 8'd47; b = 8'd2;  #10 
a = 8'd47; b = 8'd3;  #10 
a = 8'd47; b = 8'd4;  #10 
a = 8'd47; b = 8'd5;  #10 
a = 8'd47; b = 8'd6;  #10 
a = 8'd47; b = 8'd7;  #10 
a = 8'd47; b = 8'd8;  #10 
a = 8'd47; b = 8'd9;  #10 
a = 8'd47; b = 8'd10;  #10 
a = 8'd47; b = 8'd11;  #10 
a = 8'd47; b = 8'd12;  #10 
a = 8'd47; b = 8'd13;  #10 
a = 8'd47; b = 8'd14;  #10 
a = 8'd47; b = 8'd15;  #10 
a = 8'd47; b = 8'd16;  #10 
a = 8'd47; b = 8'd17;  #10 
a = 8'd47; b = 8'd18;  #10 
a = 8'd47; b = 8'd19;  #10 
a = 8'd47; b = 8'd20;  #10 
a = 8'd47; b = 8'd21;  #10 
a = 8'd47; b = 8'd22;  #10 
a = 8'd47; b = 8'd23;  #10 
a = 8'd47; b = 8'd24;  #10 
a = 8'd47; b = 8'd25;  #10 
a = 8'd47; b = 8'd26;  #10 
a = 8'd47; b = 8'd27;  #10 
a = 8'd47; b = 8'd28;  #10 
a = 8'd47; b = 8'd29;  #10 
a = 8'd47; b = 8'd30;  #10 
a = 8'd47; b = 8'd31;  #10 
a = 8'd47; b = 8'd32;  #10 
a = 8'd47; b = 8'd33;  #10 
a = 8'd47; b = 8'd34;  #10 
a = 8'd47; b = 8'd35;  #10 
a = 8'd47; b = 8'd36;  #10 
a = 8'd47; b = 8'd37;  #10 
a = 8'd47; b = 8'd38;  #10 
a = 8'd47; b = 8'd39;  #10 
a = 8'd47; b = 8'd40;  #10 
a = 8'd47; b = 8'd41;  #10 
a = 8'd47; b = 8'd42;  #10 
a = 8'd47; b = 8'd43;  #10 
a = 8'd47; b = 8'd44;  #10 
a = 8'd47; b = 8'd45;  #10 
a = 8'd47; b = 8'd46;  #10 
a = 8'd47; b = 8'd47;  #10 
a = 8'd47; b = 8'd48;  #10 
a = 8'd47; b = 8'd49;  #10 
a = 8'd47; b = 8'd50;  #10 
a = 8'd47; b = 8'd51;  #10 
a = 8'd47; b = 8'd52;  #10 
a = 8'd47; b = 8'd53;  #10 
a = 8'd47; b = 8'd54;  #10 
a = 8'd47; b = 8'd55;  #10 
a = 8'd47; b = 8'd56;  #10 
a = 8'd47; b = 8'd57;  #10 
a = 8'd47; b = 8'd58;  #10 
a = 8'd47; b = 8'd59;  #10 
a = 8'd47; b = 8'd60;  #10 
a = 8'd47; b = 8'd61;  #10 
a = 8'd47; b = 8'd62;  #10 
a = 8'd47; b = 8'd63;  #10 
a = 8'd47; b = 8'd64;  #10 
a = 8'd47; b = 8'd65;  #10 
a = 8'd47; b = 8'd66;  #10 
a = 8'd47; b = 8'd67;  #10 
a = 8'd47; b = 8'd68;  #10 
a = 8'd47; b = 8'd69;  #10 
a = 8'd47; b = 8'd70;  #10 
a = 8'd47; b = 8'd71;  #10 
a = 8'd47; b = 8'd72;  #10 
a = 8'd47; b = 8'd73;  #10 
a = 8'd47; b = 8'd74;  #10 
a = 8'd47; b = 8'd75;  #10 
a = 8'd47; b = 8'd76;  #10 
a = 8'd47; b = 8'd77;  #10 
a = 8'd47; b = 8'd78;  #10 
a = 8'd47; b = 8'd79;  #10 
a = 8'd47; b = 8'd80;  #10 
a = 8'd47; b = 8'd81;  #10 
a = 8'd47; b = 8'd82;  #10 
a = 8'd47; b = 8'd83;  #10 
a = 8'd47; b = 8'd84;  #10 
a = 8'd47; b = 8'd85;  #10 
a = 8'd47; b = 8'd86;  #10 
a = 8'd47; b = 8'd87;  #10 
a = 8'd47; b = 8'd88;  #10 
a = 8'd47; b = 8'd89;  #10 
a = 8'd47; b = 8'd90;  #10 
a = 8'd47; b = 8'd91;  #10 
a = 8'd47; b = 8'd92;  #10 
a = 8'd47; b = 8'd93;  #10 
a = 8'd47; b = 8'd94;  #10 
a = 8'd47; b = 8'd95;  #10 
a = 8'd47; b = 8'd96;  #10 
a = 8'd47; b = 8'd97;  #10 
a = 8'd47; b = 8'd98;  #10 
a = 8'd47; b = 8'd99;  #10 
a = 8'd47; b = 8'd100;  #10 
a = 8'd47; b = 8'd101;  #10 
a = 8'd47; b = 8'd102;  #10 
a = 8'd47; b = 8'd103;  #10 
a = 8'd47; b = 8'd104;  #10 
a = 8'd47; b = 8'd105;  #10 
a = 8'd47; b = 8'd106;  #10 
a = 8'd47; b = 8'd107;  #10 
a = 8'd47; b = 8'd108;  #10 
a = 8'd47; b = 8'd109;  #10 
a = 8'd47; b = 8'd110;  #10 
a = 8'd47; b = 8'd111;  #10 
a = 8'd47; b = 8'd112;  #10 
a = 8'd47; b = 8'd113;  #10 
a = 8'd47; b = 8'd114;  #10 
a = 8'd47; b = 8'd115;  #10 
a = 8'd47; b = 8'd116;  #10 
a = 8'd47; b = 8'd117;  #10 
a = 8'd47; b = 8'd118;  #10 
a = 8'd47; b = 8'd119;  #10 
a = 8'd47; b = 8'd120;  #10 
a = 8'd47; b = 8'd121;  #10 
a = 8'd47; b = 8'd122;  #10 
a = 8'd47; b = 8'd123;  #10 
a = 8'd47; b = 8'd124;  #10 
a = 8'd47; b = 8'd125;  #10 
a = 8'd47; b = 8'd126;  #10 
a = 8'd47; b = 8'd127;  #10 
a = 8'd47; b = 8'd128;  #10 
a = 8'd47; b = 8'd129;  #10 
a = 8'd47; b = 8'd130;  #10 
a = 8'd47; b = 8'd131;  #10 
a = 8'd47; b = 8'd132;  #10 
a = 8'd47; b = 8'd133;  #10 
a = 8'd47; b = 8'd134;  #10 
a = 8'd47; b = 8'd135;  #10 
a = 8'd47; b = 8'd136;  #10 
a = 8'd47; b = 8'd137;  #10 
a = 8'd47; b = 8'd138;  #10 
a = 8'd47; b = 8'd139;  #10 
a = 8'd47; b = 8'd140;  #10 
a = 8'd47; b = 8'd141;  #10 
a = 8'd47; b = 8'd142;  #10 
a = 8'd47; b = 8'd143;  #10 
a = 8'd47; b = 8'd144;  #10 
a = 8'd47; b = 8'd145;  #10 
a = 8'd47; b = 8'd146;  #10 
a = 8'd47; b = 8'd147;  #10 
a = 8'd47; b = 8'd148;  #10 
a = 8'd47; b = 8'd149;  #10 
a = 8'd47; b = 8'd150;  #10 
a = 8'd47; b = 8'd151;  #10 
a = 8'd47; b = 8'd152;  #10 
a = 8'd47; b = 8'd153;  #10 
a = 8'd47; b = 8'd154;  #10 
a = 8'd47; b = 8'd155;  #10 
a = 8'd47; b = 8'd156;  #10 
a = 8'd47; b = 8'd157;  #10 
a = 8'd47; b = 8'd158;  #10 
a = 8'd47; b = 8'd159;  #10 
a = 8'd47; b = 8'd160;  #10 
a = 8'd47; b = 8'd161;  #10 
a = 8'd47; b = 8'd162;  #10 
a = 8'd47; b = 8'd163;  #10 
a = 8'd47; b = 8'd164;  #10 
a = 8'd47; b = 8'd165;  #10 
a = 8'd47; b = 8'd166;  #10 
a = 8'd47; b = 8'd167;  #10 
a = 8'd47; b = 8'd168;  #10 
a = 8'd47; b = 8'd169;  #10 
a = 8'd47; b = 8'd170;  #10 
a = 8'd47; b = 8'd171;  #10 
a = 8'd47; b = 8'd172;  #10 
a = 8'd47; b = 8'd173;  #10 
a = 8'd47; b = 8'd174;  #10 
a = 8'd47; b = 8'd175;  #10 
a = 8'd47; b = 8'd176;  #10 
a = 8'd47; b = 8'd177;  #10 
a = 8'd47; b = 8'd178;  #10 
a = 8'd47; b = 8'd179;  #10 
a = 8'd47; b = 8'd180;  #10 
a = 8'd47; b = 8'd181;  #10 
a = 8'd47; b = 8'd182;  #10 
a = 8'd47; b = 8'd183;  #10 
a = 8'd47; b = 8'd184;  #10 
a = 8'd47; b = 8'd185;  #10 
a = 8'd47; b = 8'd186;  #10 
a = 8'd47; b = 8'd187;  #10 
a = 8'd47; b = 8'd188;  #10 
a = 8'd47; b = 8'd189;  #10 
a = 8'd47; b = 8'd190;  #10 
a = 8'd47; b = 8'd191;  #10 
a = 8'd47; b = 8'd192;  #10 
a = 8'd47; b = 8'd193;  #10 
a = 8'd47; b = 8'd194;  #10 
a = 8'd47; b = 8'd195;  #10 
a = 8'd47; b = 8'd196;  #10 
a = 8'd47; b = 8'd197;  #10 
a = 8'd47; b = 8'd198;  #10 
a = 8'd47; b = 8'd199;  #10 
a = 8'd47; b = 8'd200;  #10 
a = 8'd47; b = 8'd201;  #10 
a = 8'd47; b = 8'd202;  #10 
a = 8'd47; b = 8'd203;  #10 
a = 8'd47; b = 8'd204;  #10 
a = 8'd47; b = 8'd205;  #10 
a = 8'd47; b = 8'd206;  #10 
a = 8'd47; b = 8'd207;  #10 
a = 8'd47; b = 8'd208;  #10 
a = 8'd47; b = 8'd209;  #10 
a = 8'd47; b = 8'd210;  #10 
a = 8'd47; b = 8'd211;  #10 
a = 8'd47; b = 8'd212;  #10 
a = 8'd47; b = 8'd213;  #10 
a = 8'd47; b = 8'd214;  #10 
a = 8'd47; b = 8'd215;  #10 
a = 8'd47; b = 8'd216;  #10 
a = 8'd47; b = 8'd217;  #10 
a = 8'd47; b = 8'd218;  #10 
a = 8'd47; b = 8'd219;  #10 
a = 8'd47; b = 8'd220;  #10 
a = 8'd47; b = 8'd221;  #10 
a = 8'd47; b = 8'd222;  #10 
a = 8'd47; b = 8'd223;  #10 
a = 8'd47; b = 8'd224;  #10 
a = 8'd47; b = 8'd225;  #10 
a = 8'd47; b = 8'd226;  #10 
a = 8'd47; b = 8'd227;  #10 
a = 8'd47; b = 8'd228;  #10 
a = 8'd47; b = 8'd229;  #10 
a = 8'd47; b = 8'd230;  #10 
a = 8'd47; b = 8'd231;  #10 
a = 8'd47; b = 8'd232;  #10 
a = 8'd47; b = 8'd233;  #10 
a = 8'd47; b = 8'd234;  #10 
a = 8'd47; b = 8'd235;  #10 
a = 8'd47; b = 8'd236;  #10 
a = 8'd47; b = 8'd237;  #10 
a = 8'd47; b = 8'd238;  #10 
a = 8'd47; b = 8'd239;  #10 
a = 8'd47; b = 8'd240;  #10 
a = 8'd47; b = 8'd241;  #10 
a = 8'd47; b = 8'd242;  #10 
a = 8'd47; b = 8'd243;  #10 
a = 8'd47; b = 8'd244;  #10 
a = 8'd47; b = 8'd245;  #10 
a = 8'd47; b = 8'd246;  #10 
a = 8'd47; b = 8'd247;  #10 
a = 8'd47; b = 8'd248;  #10 
a = 8'd47; b = 8'd249;  #10 
a = 8'd47; b = 8'd250;  #10 
a = 8'd47; b = 8'd251;  #10 
a = 8'd47; b = 8'd252;  #10 
a = 8'd47; b = 8'd253;  #10 
a = 8'd47; b = 8'd254;  #10 
a = 8'd47; b = 8'd255;  #10 
a = 8'd48; b = 8'd0;  #10 
a = 8'd48; b = 8'd1;  #10 
a = 8'd48; b = 8'd2;  #10 
a = 8'd48; b = 8'd3;  #10 
a = 8'd48; b = 8'd4;  #10 
a = 8'd48; b = 8'd5;  #10 
a = 8'd48; b = 8'd6;  #10 
a = 8'd48; b = 8'd7;  #10 
a = 8'd48; b = 8'd8;  #10 
a = 8'd48; b = 8'd9;  #10 
a = 8'd48; b = 8'd10;  #10 
a = 8'd48; b = 8'd11;  #10 
a = 8'd48; b = 8'd12;  #10 
a = 8'd48; b = 8'd13;  #10 
a = 8'd48; b = 8'd14;  #10 
a = 8'd48; b = 8'd15;  #10 
a = 8'd48; b = 8'd16;  #10 
a = 8'd48; b = 8'd17;  #10 
a = 8'd48; b = 8'd18;  #10 
a = 8'd48; b = 8'd19;  #10 
a = 8'd48; b = 8'd20;  #10 
a = 8'd48; b = 8'd21;  #10 
a = 8'd48; b = 8'd22;  #10 
a = 8'd48; b = 8'd23;  #10 
a = 8'd48; b = 8'd24;  #10 
a = 8'd48; b = 8'd25;  #10 
a = 8'd48; b = 8'd26;  #10 
a = 8'd48; b = 8'd27;  #10 
a = 8'd48; b = 8'd28;  #10 
a = 8'd48; b = 8'd29;  #10 
a = 8'd48; b = 8'd30;  #10 
a = 8'd48; b = 8'd31;  #10 
a = 8'd48; b = 8'd32;  #10 
a = 8'd48; b = 8'd33;  #10 
a = 8'd48; b = 8'd34;  #10 
a = 8'd48; b = 8'd35;  #10 
a = 8'd48; b = 8'd36;  #10 
a = 8'd48; b = 8'd37;  #10 
a = 8'd48; b = 8'd38;  #10 
a = 8'd48; b = 8'd39;  #10 
a = 8'd48; b = 8'd40;  #10 
a = 8'd48; b = 8'd41;  #10 
a = 8'd48; b = 8'd42;  #10 
a = 8'd48; b = 8'd43;  #10 
a = 8'd48; b = 8'd44;  #10 
a = 8'd48; b = 8'd45;  #10 
a = 8'd48; b = 8'd46;  #10 
a = 8'd48; b = 8'd47;  #10 
a = 8'd48; b = 8'd48;  #10 
a = 8'd48; b = 8'd49;  #10 
a = 8'd48; b = 8'd50;  #10 
a = 8'd48; b = 8'd51;  #10 
a = 8'd48; b = 8'd52;  #10 
a = 8'd48; b = 8'd53;  #10 
a = 8'd48; b = 8'd54;  #10 
a = 8'd48; b = 8'd55;  #10 
a = 8'd48; b = 8'd56;  #10 
a = 8'd48; b = 8'd57;  #10 
a = 8'd48; b = 8'd58;  #10 
a = 8'd48; b = 8'd59;  #10 
a = 8'd48; b = 8'd60;  #10 
a = 8'd48; b = 8'd61;  #10 
a = 8'd48; b = 8'd62;  #10 
a = 8'd48; b = 8'd63;  #10 
a = 8'd48; b = 8'd64;  #10 
a = 8'd48; b = 8'd65;  #10 
a = 8'd48; b = 8'd66;  #10 
a = 8'd48; b = 8'd67;  #10 
a = 8'd48; b = 8'd68;  #10 
a = 8'd48; b = 8'd69;  #10 
a = 8'd48; b = 8'd70;  #10 
a = 8'd48; b = 8'd71;  #10 
a = 8'd48; b = 8'd72;  #10 
a = 8'd48; b = 8'd73;  #10 
a = 8'd48; b = 8'd74;  #10 
a = 8'd48; b = 8'd75;  #10 
a = 8'd48; b = 8'd76;  #10 
a = 8'd48; b = 8'd77;  #10 
a = 8'd48; b = 8'd78;  #10 
a = 8'd48; b = 8'd79;  #10 
a = 8'd48; b = 8'd80;  #10 
a = 8'd48; b = 8'd81;  #10 
a = 8'd48; b = 8'd82;  #10 
a = 8'd48; b = 8'd83;  #10 
a = 8'd48; b = 8'd84;  #10 
a = 8'd48; b = 8'd85;  #10 
a = 8'd48; b = 8'd86;  #10 
a = 8'd48; b = 8'd87;  #10 
a = 8'd48; b = 8'd88;  #10 
a = 8'd48; b = 8'd89;  #10 
a = 8'd48; b = 8'd90;  #10 
a = 8'd48; b = 8'd91;  #10 
a = 8'd48; b = 8'd92;  #10 
a = 8'd48; b = 8'd93;  #10 
a = 8'd48; b = 8'd94;  #10 
a = 8'd48; b = 8'd95;  #10 
a = 8'd48; b = 8'd96;  #10 
a = 8'd48; b = 8'd97;  #10 
a = 8'd48; b = 8'd98;  #10 
a = 8'd48; b = 8'd99;  #10 
a = 8'd48; b = 8'd100;  #10 
a = 8'd48; b = 8'd101;  #10 
a = 8'd48; b = 8'd102;  #10 
a = 8'd48; b = 8'd103;  #10 
a = 8'd48; b = 8'd104;  #10 
a = 8'd48; b = 8'd105;  #10 
a = 8'd48; b = 8'd106;  #10 
a = 8'd48; b = 8'd107;  #10 
a = 8'd48; b = 8'd108;  #10 
a = 8'd48; b = 8'd109;  #10 
a = 8'd48; b = 8'd110;  #10 
a = 8'd48; b = 8'd111;  #10 
a = 8'd48; b = 8'd112;  #10 
a = 8'd48; b = 8'd113;  #10 
a = 8'd48; b = 8'd114;  #10 
a = 8'd48; b = 8'd115;  #10 
a = 8'd48; b = 8'd116;  #10 
a = 8'd48; b = 8'd117;  #10 
a = 8'd48; b = 8'd118;  #10 
a = 8'd48; b = 8'd119;  #10 
a = 8'd48; b = 8'd120;  #10 
a = 8'd48; b = 8'd121;  #10 
a = 8'd48; b = 8'd122;  #10 
a = 8'd48; b = 8'd123;  #10 
a = 8'd48; b = 8'd124;  #10 
a = 8'd48; b = 8'd125;  #10 
a = 8'd48; b = 8'd126;  #10 
a = 8'd48; b = 8'd127;  #10 
a = 8'd48; b = 8'd128;  #10 
a = 8'd48; b = 8'd129;  #10 
a = 8'd48; b = 8'd130;  #10 
a = 8'd48; b = 8'd131;  #10 
a = 8'd48; b = 8'd132;  #10 
a = 8'd48; b = 8'd133;  #10 
a = 8'd48; b = 8'd134;  #10 
a = 8'd48; b = 8'd135;  #10 
a = 8'd48; b = 8'd136;  #10 
a = 8'd48; b = 8'd137;  #10 
a = 8'd48; b = 8'd138;  #10 
a = 8'd48; b = 8'd139;  #10 
a = 8'd48; b = 8'd140;  #10 
a = 8'd48; b = 8'd141;  #10 
a = 8'd48; b = 8'd142;  #10 
a = 8'd48; b = 8'd143;  #10 
a = 8'd48; b = 8'd144;  #10 
a = 8'd48; b = 8'd145;  #10 
a = 8'd48; b = 8'd146;  #10 
a = 8'd48; b = 8'd147;  #10 
a = 8'd48; b = 8'd148;  #10 
a = 8'd48; b = 8'd149;  #10 
a = 8'd48; b = 8'd150;  #10 
a = 8'd48; b = 8'd151;  #10 
a = 8'd48; b = 8'd152;  #10 
a = 8'd48; b = 8'd153;  #10 
a = 8'd48; b = 8'd154;  #10 
a = 8'd48; b = 8'd155;  #10 
a = 8'd48; b = 8'd156;  #10 
a = 8'd48; b = 8'd157;  #10 
a = 8'd48; b = 8'd158;  #10 
a = 8'd48; b = 8'd159;  #10 
a = 8'd48; b = 8'd160;  #10 
a = 8'd48; b = 8'd161;  #10 
a = 8'd48; b = 8'd162;  #10 
a = 8'd48; b = 8'd163;  #10 
a = 8'd48; b = 8'd164;  #10 
a = 8'd48; b = 8'd165;  #10 
a = 8'd48; b = 8'd166;  #10 
a = 8'd48; b = 8'd167;  #10 
a = 8'd48; b = 8'd168;  #10 
a = 8'd48; b = 8'd169;  #10 
a = 8'd48; b = 8'd170;  #10 
a = 8'd48; b = 8'd171;  #10 
a = 8'd48; b = 8'd172;  #10 
a = 8'd48; b = 8'd173;  #10 
a = 8'd48; b = 8'd174;  #10 
a = 8'd48; b = 8'd175;  #10 
a = 8'd48; b = 8'd176;  #10 
a = 8'd48; b = 8'd177;  #10 
a = 8'd48; b = 8'd178;  #10 
a = 8'd48; b = 8'd179;  #10 
a = 8'd48; b = 8'd180;  #10 
a = 8'd48; b = 8'd181;  #10 
a = 8'd48; b = 8'd182;  #10 
a = 8'd48; b = 8'd183;  #10 
a = 8'd48; b = 8'd184;  #10 
a = 8'd48; b = 8'd185;  #10 
a = 8'd48; b = 8'd186;  #10 
a = 8'd48; b = 8'd187;  #10 
a = 8'd48; b = 8'd188;  #10 
a = 8'd48; b = 8'd189;  #10 
a = 8'd48; b = 8'd190;  #10 
a = 8'd48; b = 8'd191;  #10 
a = 8'd48; b = 8'd192;  #10 
a = 8'd48; b = 8'd193;  #10 
a = 8'd48; b = 8'd194;  #10 
a = 8'd48; b = 8'd195;  #10 
a = 8'd48; b = 8'd196;  #10 
a = 8'd48; b = 8'd197;  #10 
a = 8'd48; b = 8'd198;  #10 
a = 8'd48; b = 8'd199;  #10 
a = 8'd48; b = 8'd200;  #10 
a = 8'd48; b = 8'd201;  #10 
a = 8'd48; b = 8'd202;  #10 
a = 8'd48; b = 8'd203;  #10 
a = 8'd48; b = 8'd204;  #10 
a = 8'd48; b = 8'd205;  #10 
a = 8'd48; b = 8'd206;  #10 
a = 8'd48; b = 8'd207;  #10 
a = 8'd48; b = 8'd208;  #10 
a = 8'd48; b = 8'd209;  #10 
a = 8'd48; b = 8'd210;  #10 
a = 8'd48; b = 8'd211;  #10 
a = 8'd48; b = 8'd212;  #10 
a = 8'd48; b = 8'd213;  #10 
a = 8'd48; b = 8'd214;  #10 
a = 8'd48; b = 8'd215;  #10 
a = 8'd48; b = 8'd216;  #10 
a = 8'd48; b = 8'd217;  #10 
a = 8'd48; b = 8'd218;  #10 
a = 8'd48; b = 8'd219;  #10 
a = 8'd48; b = 8'd220;  #10 
a = 8'd48; b = 8'd221;  #10 
a = 8'd48; b = 8'd222;  #10 
a = 8'd48; b = 8'd223;  #10 
a = 8'd48; b = 8'd224;  #10 
a = 8'd48; b = 8'd225;  #10 
a = 8'd48; b = 8'd226;  #10 
a = 8'd48; b = 8'd227;  #10 
a = 8'd48; b = 8'd228;  #10 
a = 8'd48; b = 8'd229;  #10 
a = 8'd48; b = 8'd230;  #10 
a = 8'd48; b = 8'd231;  #10 
a = 8'd48; b = 8'd232;  #10 
a = 8'd48; b = 8'd233;  #10 
a = 8'd48; b = 8'd234;  #10 
a = 8'd48; b = 8'd235;  #10 
a = 8'd48; b = 8'd236;  #10 
a = 8'd48; b = 8'd237;  #10 
a = 8'd48; b = 8'd238;  #10 
a = 8'd48; b = 8'd239;  #10 
a = 8'd48; b = 8'd240;  #10 
a = 8'd48; b = 8'd241;  #10 
a = 8'd48; b = 8'd242;  #10 
a = 8'd48; b = 8'd243;  #10 
a = 8'd48; b = 8'd244;  #10 
a = 8'd48; b = 8'd245;  #10 
a = 8'd48; b = 8'd246;  #10 
a = 8'd48; b = 8'd247;  #10 
a = 8'd48; b = 8'd248;  #10 
a = 8'd48; b = 8'd249;  #10 
a = 8'd48; b = 8'd250;  #10 
a = 8'd48; b = 8'd251;  #10 
a = 8'd48; b = 8'd252;  #10 
a = 8'd48; b = 8'd253;  #10 
a = 8'd48; b = 8'd254;  #10 
a = 8'd48; b = 8'd255;  #10 
a = 8'd49; b = 8'd0;  #10 
a = 8'd49; b = 8'd1;  #10 
a = 8'd49; b = 8'd2;  #10 
a = 8'd49; b = 8'd3;  #10 
a = 8'd49; b = 8'd4;  #10 
a = 8'd49; b = 8'd5;  #10 
a = 8'd49; b = 8'd6;  #10 
a = 8'd49; b = 8'd7;  #10 
a = 8'd49; b = 8'd8;  #10 
a = 8'd49; b = 8'd9;  #10 
a = 8'd49; b = 8'd10;  #10 
a = 8'd49; b = 8'd11;  #10 
a = 8'd49; b = 8'd12;  #10 
a = 8'd49; b = 8'd13;  #10 
a = 8'd49; b = 8'd14;  #10 
a = 8'd49; b = 8'd15;  #10 
a = 8'd49; b = 8'd16;  #10 
a = 8'd49; b = 8'd17;  #10 
a = 8'd49; b = 8'd18;  #10 
a = 8'd49; b = 8'd19;  #10 
a = 8'd49; b = 8'd20;  #10 
a = 8'd49; b = 8'd21;  #10 
a = 8'd49; b = 8'd22;  #10 
a = 8'd49; b = 8'd23;  #10 
a = 8'd49; b = 8'd24;  #10 
a = 8'd49; b = 8'd25;  #10 
a = 8'd49; b = 8'd26;  #10 
a = 8'd49; b = 8'd27;  #10 
a = 8'd49; b = 8'd28;  #10 
a = 8'd49; b = 8'd29;  #10 
a = 8'd49; b = 8'd30;  #10 
a = 8'd49; b = 8'd31;  #10 
a = 8'd49; b = 8'd32;  #10 
a = 8'd49; b = 8'd33;  #10 
a = 8'd49; b = 8'd34;  #10 
a = 8'd49; b = 8'd35;  #10 
a = 8'd49; b = 8'd36;  #10 
a = 8'd49; b = 8'd37;  #10 
a = 8'd49; b = 8'd38;  #10 
a = 8'd49; b = 8'd39;  #10 
a = 8'd49; b = 8'd40;  #10 
a = 8'd49; b = 8'd41;  #10 
a = 8'd49; b = 8'd42;  #10 
a = 8'd49; b = 8'd43;  #10 
a = 8'd49; b = 8'd44;  #10 
a = 8'd49; b = 8'd45;  #10 
a = 8'd49; b = 8'd46;  #10 
a = 8'd49; b = 8'd47;  #10 
a = 8'd49; b = 8'd48;  #10 
a = 8'd49; b = 8'd49;  #10 
a = 8'd49; b = 8'd50;  #10 
a = 8'd49; b = 8'd51;  #10 
a = 8'd49; b = 8'd52;  #10 
a = 8'd49; b = 8'd53;  #10 
a = 8'd49; b = 8'd54;  #10 
a = 8'd49; b = 8'd55;  #10 
a = 8'd49; b = 8'd56;  #10 
a = 8'd49; b = 8'd57;  #10 
a = 8'd49; b = 8'd58;  #10 
a = 8'd49; b = 8'd59;  #10 
a = 8'd49; b = 8'd60;  #10 
a = 8'd49; b = 8'd61;  #10 
a = 8'd49; b = 8'd62;  #10 
a = 8'd49; b = 8'd63;  #10 
a = 8'd49; b = 8'd64;  #10 
a = 8'd49; b = 8'd65;  #10 
a = 8'd49; b = 8'd66;  #10 
a = 8'd49; b = 8'd67;  #10 
a = 8'd49; b = 8'd68;  #10 
a = 8'd49; b = 8'd69;  #10 
a = 8'd49; b = 8'd70;  #10 
a = 8'd49; b = 8'd71;  #10 
a = 8'd49; b = 8'd72;  #10 
a = 8'd49; b = 8'd73;  #10 
a = 8'd49; b = 8'd74;  #10 
a = 8'd49; b = 8'd75;  #10 
a = 8'd49; b = 8'd76;  #10 
a = 8'd49; b = 8'd77;  #10 
a = 8'd49; b = 8'd78;  #10 
a = 8'd49; b = 8'd79;  #10 
a = 8'd49; b = 8'd80;  #10 
a = 8'd49; b = 8'd81;  #10 
a = 8'd49; b = 8'd82;  #10 
a = 8'd49; b = 8'd83;  #10 
a = 8'd49; b = 8'd84;  #10 
a = 8'd49; b = 8'd85;  #10 
a = 8'd49; b = 8'd86;  #10 
a = 8'd49; b = 8'd87;  #10 
a = 8'd49; b = 8'd88;  #10 
a = 8'd49; b = 8'd89;  #10 
a = 8'd49; b = 8'd90;  #10 
a = 8'd49; b = 8'd91;  #10 
a = 8'd49; b = 8'd92;  #10 
a = 8'd49; b = 8'd93;  #10 
a = 8'd49; b = 8'd94;  #10 
a = 8'd49; b = 8'd95;  #10 
a = 8'd49; b = 8'd96;  #10 
a = 8'd49; b = 8'd97;  #10 
a = 8'd49; b = 8'd98;  #10 
a = 8'd49; b = 8'd99;  #10 
a = 8'd49; b = 8'd100;  #10 
a = 8'd49; b = 8'd101;  #10 
a = 8'd49; b = 8'd102;  #10 
a = 8'd49; b = 8'd103;  #10 
a = 8'd49; b = 8'd104;  #10 
a = 8'd49; b = 8'd105;  #10 
a = 8'd49; b = 8'd106;  #10 
a = 8'd49; b = 8'd107;  #10 
a = 8'd49; b = 8'd108;  #10 
a = 8'd49; b = 8'd109;  #10 
a = 8'd49; b = 8'd110;  #10 
a = 8'd49; b = 8'd111;  #10 
a = 8'd49; b = 8'd112;  #10 
a = 8'd49; b = 8'd113;  #10 
a = 8'd49; b = 8'd114;  #10 
a = 8'd49; b = 8'd115;  #10 
a = 8'd49; b = 8'd116;  #10 
a = 8'd49; b = 8'd117;  #10 
a = 8'd49; b = 8'd118;  #10 
a = 8'd49; b = 8'd119;  #10 
a = 8'd49; b = 8'd120;  #10 
a = 8'd49; b = 8'd121;  #10 
a = 8'd49; b = 8'd122;  #10 
a = 8'd49; b = 8'd123;  #10 
a = 8'd49; b = 8'd124;  #10 
a = 8'd49; b = 8'd125;  #10 
a = 8'd49; b = 8'd126;  #10 
a = 8'd49; b = 8'd127;  #10 
a = 8'd49; b = 8'd128;  #10 
a = 8'd49; b = 8'd129;  #10 
a = 8'd49; b = 8'd130;  #10 
a = 8'd49; b = 8'd131;  #10 
a = 8'd49; b = 8'd132;  #10 
a = 8'd49; b = 8'd133;  #10 
a = 8'd49; b = 8'd134;  #10 
a = 8'd49; b = 8'd135;  #10 
a = 8'd49; b = 8'd136;  #10 
a = 8'd49; b = 8'd137;  #10 
a = 8'd49; b = 8'd138;  #10 
a = 8'd49; b = 8'd139;  #10 
a = 8'd49; b = 8'd140;  #10 
a = 8'd49; b = 8'd141;  #10 
a = 8'd49; b = 8'd142;  #10 
a = 8'd49; b = 8'd143;  #10 
a = 8'd49; b = 8'd144;  #10 
a = 8'd49; b = 8'd145;  #10 
a = 8'd49; b = 8'd146;  #10 
a = 8'd49; b = 8'd147;  #10 
a = 8'd49; b = 8'd148;  #10 
a = 8'd49; b = 8'd149;  #10 
a = 8'd49; b = 8'd150;  #10 
a = 8'd49; b = 8'd151;  #10 
a = 8'd49; b = 8'd152;  #10 
a = 8'd49; b = 8'd153;  #10 
a = 8'd49; b = 8'd154;  #10 
a = 8'd49; b = 8'd155;  #10 
a = 8'd49; b = 8'd156;  #10 
a = 8'd49; b = 8'd157;  #10 
a = 8'd49; b = 8'd158;  #10 
a = 8'd49; b = 8'd159;  #10 
a = 8'd49; b = 8'd160;  #10 
a = 8'd49; b = 8'd161;  #10 
a = 8'd49; b = 8'd162;  #10 
a = 8'd49; b = 8'd163;  #10 
a = 8'd49; b = 8'd164;  #10 
a = 8'd49; b = 8'd165;  #10 
a = 8'd49; b = 8'd166;  #10 
a = 8'd49; b = 8'd167;  #10 
a = 8'd49; b = 8'd168;  #10 
a = 8'd49; b = 8'd169;  #10 
a = 8'd49; b = 8'd170;  #10 
a = 8'd49; b = 8'd171;  #10 
a = 8'd49; b = 8'd172;  #10 
a = 8'd49; b = 8'd173;  #10 
a = 8'd49; b = 8'd174;  #10 
a = 8'd49; b = 8'd175;  #10 
a = 8'd49; b = 8'd176;  #10 
a = 8'd49; b = 8'd177;  #10 
a = 8'd49; b = 8'd178;  #10 
a = 8'd49; b = 8'd179;  #10 
a = 8'd49; b = 8'd180;  #10 
a = 8'd49; b = 8'd181;  #10 
a = 8'd49; b = 8'd182;  #10 
a = 8'd49; b = 8'd183;  #10 
a = 8'd49; b = 8'd184;  #10 
a = 8'd49; b = 8'd185;  #10 
a = 8'd49; b = 8'd186;  #10 
a = 8'd49; b = 8'd187;  #10 
a = 8'd49; b = 8'd188;  #10 
a = 8'd49; b = 8'd189;  #10 
a = 8'd49; b = 8'd190;  #10 
a = 8'd49; b = 8'd191;  #10 
a = 8'd49; b = 8'd192;  #10 
a = 8'd49; b = 8'd193;  #10 
a = 8'd49; b = 8'd194;  #10 
a = 8'd49; b = 8'd195;  #10 
a = 8'd49; b = 8'd196;  #10 
a = 8'd49; b = 8'd197;  #10 
a = 8'd49; b = 8'd198;  #10 
a = 8'd49; b = 8'd199;  #10 
a = 8'd49; b = 8'd200;  #10 
a = 8'd49; b = 8'd201;  #10 
a = 8'd49; b = 8'd202;  #10 
a = 8'd49; b = 8'd203;  #10 
a = 8'd49; b = 8'd204;  #10 
a = 8'd49; b = 8'd205;  #10 
a = 8'd49; b = 8'd206;  #10 
a = 8'd49; b = 8'd207;  #10 
a = 8'd49; b = 8'd208;  #10 
a = 8'd49; b = 8'd209;  #10 
a = 8'd49; b = 8'd210;  #10 
a = 8'd49; b = 8'd211;  #10 
a = 8'd49; b = 8'd212;  #10 
a = 8'd49; b = 8'd213;  #10 
a = 8'd49; b = 8'd214;  #10 
a = 8'd49; b = 8'd215;  #10 
a = 8'd49; b = 8'd216;  #10 
a = 8'd49; b = 8'd217;  #10 
a = 8'd49; b = 8'd218;  #10 
a = 8'd49; b = 8'd219;  #10 
a = 8'd49; b = 8'd220;  #10 
a = 8'd49; b = 8'd221;  #10 
a = 8'd49; b = 8'd222;  #10 
a = 8'd49; b = 8'd223;  #10 
a = 8'd49; b = 8'd224;  #10 
a = 8'd49; b = 8'd225;  #10 
a = 8'd49; b = 8'd226;  #10 
a = 8'd49; b = 8'd227;  #10 
a = 8'd49; b = 8'd228;  #10 
a = 8'd49; b = 8'd229;  #10 
a = 8'd49; b = 8'd230;  #10 
a = 8'd49; b = 8'd231;  #10 
a = 8'd49; b = 8'd232;  #10 
a = 8'd49; b = 8'd233;  #10 
a = 8'd49; b = 8'd234;  #10 
a = 8'd49; b = 8'd235;  #10 
a = 8'd49; b = 8'd236;  #10 
a = 8'd49; b = 8'd237;  #10 
a = 8'd49; b = 8'd238;  #10 
a = 8'd49; b = 8'd239;  #10 
a = 8'd49; b = 8'd240;  #10 
a = 8'd49; b = 8'd241;  #10 
a = 8'd49; b = 8'd242;  #10 
a = 8'd49; b = 8'd243;  #10 
a = 8'd49; b = 8'd244;  #10 
a = 8'd49; b = 8'd245;  #10 
a = 8'd49; b = 8'd246;  #10 
a = 8'd49; b = 8'd247;  #10 
a = 8'd49; b = 8'd248;  #10 
a = 8'd49; b = 8'd249;  #10 
a = 8'd49; b = 8'd250;  #10 
a = 8'd49; b = 8'd251;  #10 
a = 8'd49; b = 8'd252;  #10 
a = 8'd49; b = 8'd253;  #10 
a = 8'd49; b = 8'd254;  #10 
a = 8'd49; b = 8'd255;  #10 
a = 8'd50; b = 8'd0;  #10 
a = 8'd50; b = 8'd1;  #10 
a = 8'd50; b = 8'd2;  #10 
a = 8'd50; b = 8'd3;  #10 
a = 8'd50; b = 8'd4;  #10 
a = 8'd50; b = 8'd5;  #10 
a = 8'd50; b = 8'd6;  #10 
a = 8'd50; b = 8'd7;  #10 
a = 8'd50; b = 8'd8;  #10 
a = 8'd50; b = 8'd9;  #10 
a = 8'd50; b = 8'd10;  #10 
a = 8'd50; b = 8'd11;  #10 
a = 8'd50; b = 8'd12;  #10 
a = 8'd50; b = 8'd13;  #10 
a = 8'd50; b = 8'd14;  #10 
a = 8'd50; b = 8'd15;  #10 
a = 8'd50; b = 8'd16;  #10 
a = 8'd50; b = 8'd17;  #10 
a = 8'd50; b = 8'd18;  #10 
a = 8'd50; b = 8'd19;  #10 
a = 8'd50; b = 8'd20;  #10 
a = 8'd50; b = 8'd21;  #10 
a = 8'd50; b = 8'd22;  #10 
a = 8'd50; b = 8'd23;  #10 
a = 8'd50; b = 8'd24;  #10 
a = 8'd50; b = 8'd25;  #10 
a = 8'd50; b = 8'd26;  #10 
a = 8'd50; b = 8'd27;  #10 
a = 8'd50; b = 8'd28;  #10 
a = 8'd50; b = 8'd29;  #10 
a = 8'd50; b = 8'd30;  #10 
a = 8'd50; b = 8'd31;  #10 
a = 8'd50; b = 8'd32;  #10 
a = 8'd50; b = 8'd33;  #10 
a = 8'd50; b = 8'd34;  #10 
a = 8'd50; b = 8'd35;  #10 
a = 8'd50; b = 8'd36;  #10 
a = 8'd50; b = 8'd37;  #10 
a = 8'd50; b = 8'd38;  #10 
a = 8'd50; b = 8'd39;  #10 
a = 8'd50; b = 8'd40;  #10 
a = 8'd50; b = 8'd41;  #10 
a = 8'd50; b = 8'd42;  #10 
a = 8'd50; b = 8'd43;  #10 
a = 8'd50; b = 8'd44;  #10 
a = 8'd50; b = 8'd45;  #10 
a = 8'd50; b = 8'd46;  #10 
a = 8'd50; b = 8'd47;  #10 
a = 8'd50; b = 8'd48;  #10 
a = 8'd50; b = 8'd49;  #10 
a = 8'd50; b = 8'd50;  #10 
a = 8'd50; b = 8'd51;  #10 
a = 8'd50; b = 8'd52;  #10 
a = 8'd50; b = 8'd53;  #10 
a = 8'd50; b = 8'd54;  #10 
a = 8'd50; b = 8'd55;  #10 
a = 8'd50; b = 8'd56;  #10 
a = 8'd50; b = 8'd57;  #10 
a = 8'd50; b = 8'd58;  #10 
a = 8'd50; b = 8'd59;  #10 
a = 8'd50; b = 8'd60;  #10 
a = 8'd50; b = 8'd61;  #10 
a = 8'd50; b = 8'd62;  #10 
a = 8'd50; b = 8'd63;  #10 
a = 8'd50; b = 8'd64;  #10 
a = 8'd50; b = 8'd65;  #10 
a = 8'd50; b = 8'd66;  #10 
a = 8'd50; b = 8'd67;  #10 
a = 8'd50; b = 8'd68;  #10 
a = 8'd50; b = 8'd69;  #10 
a = 8'd50; b = 8'd70;  #10 
a = 8'd50; b = 8'd71;  #10 
a = 8'd50; b = 8'd72;  #10 
a = 8'd50; b = 8'd73;  #10 
a = 8'd50; b = 8'd74;  #10 
a = 8'd50; b = 8'd75;  #10 
a = 8'd50; b = 8'd76;  #10 
a = 8'd50; b = 8'd77;  #10 
a = 8'd50; b = 8'd78;  #10 
a = 8'd50; b = 8'd79;  #10 
a = 8'd50; b = 8'd80;  #10 
a = 8'd50; b = 8'd81;  #10 
a = 8'd50; b = 8'd82;  #10 
a = 8'd50; b = 8'd83;  #10 
a = 8'd50; b = 8'd84;  #10 
a = 8'd50; b = 8'd85;  #10 
a = 8'd50; b = 8'd86;  #10 
a = 8'd50; b = 8'd87;  #10 
a = 8'd50; b = 8'd88;  #10 
a = 8'd50; b = 8'd89;  #10 
a = 8'd50; b = 8'd90;  #10 
a = 8'd50; b = 8'd91;  #10 
a = 8'd50; b = 8'd92;  #10 
a = 8'd50; b = 8'd93;  #10 
a = 8'd50; b = 8'd94;  #10 
a = 8'd50; b = 8'd95;  #10 
a = 8'd50; b = 8'd96;  #10 
a = 8'd50; b = 8'd97;  #10 
a = 8'd50; b = 8'd98;  #10 
a = 8'd50; b = 8'd99;  #10 
a = 8'd50; b = 8'd100;  #10 
a = 8'd50; b = 8'd101;  #10 
a = 8'd50; b = 8'd102;  #10 
a = 8'd50; b = 8'd103;  #10 
a = 8'd50; b = 8'd104;  #10 
a = 8'd50; b = 8'd105;  #10 
a = 8'd50; b = 8'd106;  #10 
a = 8'd50; b = 8'd107;  #10 
a = 8'd50; b = 8'd108;  #10 
a = 8'd50; b = 8'd109;  #10 
a = 8'd50; b = 8'd110;  #10 
a = 8'd50; b = 8'd111;  #10 
a = 8'd50; b = 8'd112;  #10 
a = 8'd50; b = 8'd113;  #10 
a = 8'd50; b = 8'd114;  #10 
a = 8'd50; b = 8'd115;  #10 
a = 8'd50; b = 8'd116;  #10 
a = 8'd50; b = 8'd117;  #10 
a = 8'd50; b = 8'd118;  #10 
a = 8'd50; b = 8'd119;  #10 
a = 8'd50; b = 8'd120;  #10 
a = 8'd50; b = 8'd121;  #10 
a = 8'd50; b = 8'd122;  #10 
a = 8'd50; b = 8'd123;  #10 
a = 8'd50; b = 8'd124;  #10 
a = 8'd50; b = 8'd125;  #10 
a = 8'd50; b = 8'd126;  #10 
a = 8'd50; b = 8'd127;  #10 
a = 8'd50; b = 8'd128;  #10 
a = 8'd50; b = 8'd129;  #10 
a = 8'd50; b = 8'd130;  #10 
a = 8'd50; b = 8'd131;  #10 
a = 8'd50; b = 8'd132;  #10 
a = 8'd50; b = 8'd133;  #10 
a = 8'd50; b = 8'd134;  #10 
a = 8'd50; b = 8'd135;  #10 
a = 8'd50; b = 8'd136;  #10 
a = 8'd50; b = 8'd137;  #10 
a = 8'd50; b = 8'd138;  #10 
a = 8'd50; b = 8'd139;  #10 
a = 8'd50; b = 8'd140;  #10 
a = 8'd50; b = 8'd141;  #10 
a = 8'd50; b = 8'd142;  #10 
a = 8'd50; b = 8'd143;  #10 
a = 8'd50; b = 8'd144;  #10 
a = 8'd50; b = 8'd145;  #10 
a = 8'd50; b = 8'd146;  #10 
a = 8'd50; b = 8'd147;  #10 
a = 8'd50; b = 8'd148;  #10 
a = 8'd50; b = 8'd149;  #10 
a = 8'd50; b = 8'd150;  #10 
a = 8'd50; b = 8'd151;  #10 
a = 8'd50; b = 8'd152;  #10 
a = 8'd50; b = 8'd153;  #10 
a = 8'd50; b = 8'd154;  #10 
a = 8'd50; b = 8'd155;  #10 
a = 8'd50; b = 8'd156;  #10 
a = 8'd50; b = 8'd157;  #10 
a = 8'd50; b = 8'd158;  #10 
a = 8'd50; b = 8'd159;  #10 
a = 8'd50; b = 8'd160;  #10 
a = 8'd50; b = 8'd161;  #10 
a = 8'd50; b = 8'd162;  #10 
a = 8'd50; b = 8'd163;  #10 
a = 8'd50; b = 8'd164;  #10 
a = 8'd50; b = 8'd165;  #10 
a = 8'd50; b = 8'd166;  #10 
a = 8'd50; b = 8'd167;  #10 
a = 8'd50; b = 8'd168;  #10 
a = 8'd50; b = 8'd169;  #10 
a = 8'd50; b = 8'd170;  #10 
a = 8'd50; b = 8'd171;  #10 
a = 8'd50; b = 8'd172;  #10 
a = 8'd50; b = 8'd173;  #10 
a = 8'd50; b = 8'd174;  #10 
a = 8'd50; b = 8'd175;  #10 
a = 8'd50; b = 8'd176;  #10 
a = 8'd50; b = 8'd177;  #10 
a = 8'd50; b = 8'd178;  #10 
a = 8'd50; b = 8'd179;  #10 
a = 8'd50; b = 8'd180;  #10 
a = 8'd50; b = 8'd181;  #10 
a = 8'd50; b = 8'd182;  #10 
a = 8'd50; b = 8'd183;  #10 
a = 8'd50; b = 8'd184;  #10 
a = 8'd50; b = 8'd185;  #10 
a = 8'd50; b = 8'd186;  #10 
a = 8'd50; b = 8'd187;  #10 
a = 8'd50; b = 8'd188;  #10 
a = 8'd50; b = 8'd189;  #10 
a = 8'd50; b = 8'd190;  #10 
a = 8'd50; b = 8'd191;  #10 
a = 8'd50; b = 8'd192;  #10 
a = 8'd50; b = 8'd193;  #10 
a = 8'd50; b = 8'd194;  #10 
a = 8'd50; b = 8'd195;  #10 
a = 8'd50; b = 8'd196;  #10 
a = 8'd50; b = 8'd197;  #10 
a = 8'd50; b = 8'd198;  #10 
a = 8'd50; b = 8'd199;  #10 
a = 8'd50; b = 8'd200;  #10 
a = 8'd50; b = 8'd201;  #10 
a = 8'd50; b = 8'd202;  #10 
a = 8'd50; b = 8'd203;  #10 
a = 8'd50; b = 8'd204;  #10 
a = 8'd50; b = 8'd205;  #10 
a = 8'd50; b = 8'd206;  #10 
a = 8'd50; b = 8'd207;  #10 
a = 8'd50; b = 8'd208;  #10 
a = 8'd50; b = 8'd209;  #10 
a = 8'd50; b = 8'd210;  #10 
a = 8'd50; b = 8'd211;  #10 
a = 8'd50; b = 8'd212;  #10 
a = 8'd50; b = 8'd213;  #10 
a = 8'd50; b = 8'd214;  #10 
a = 8'd50; b = 8'd215;  #10 
a = 8'd50; b = 8'd216;  #10 
a = 8'd50; b = 8'd217;  #10 
a = 8'd50; b = 8'd218;  #10 
a = 8'd50; b = 8'd219;  #10 
a = 8'd50; b = 8'd220;  #10 
a = 8'd50; b = 8'd221;  #10 
a = 8'd50; b = 8'd222;  #10 
a = 8'd50; b = 8'd223;  #10 
a = 8'd50; b = 8'd224;  #10 
a = 8'd50; b = 8'd225;  #10 
a = 8'd50; b = 8'd226;  #10 
a = 8'd50; b = 8'd227;  #10 
a = 8'd50; b = 8'd228;  #10 
a = 8'd50; b = 8'd229;  #10 
a = 8'd50; b = 8'd230;  #10 
a = 8'd50; b = 8'd231;  #10 
a = 8'd50; b = 8'd232;  #10 
a = 8'd50; b = 8'd233;  #10 
a = 8'd50; b = 8'd234;  #10 
a = 8'd50; b = 8'd235;  #10 
a = 8'd50; b = 8'd236;  #10 
a = 8'd50; b = 8'd237;  #10 
a = 8'd50; b = 8'd238;  #10 
a = 8'd50; b = 8'd239;  #10 
a = 8'd50; b = 8'd240;  #10 
a = 8'd50; b = 8'd241;  #10 
a = 8'd50; b = 8'd242;  #10 
a = 8'd50; b = 8'd243;  #10 
a = 8'd50; b = 8'd244;  #10 
a = 8'd50; b = 8'd245;  #10 
a = 8'd50; b = 8'd246;  #10 
a = 8'd50; b = 8'd247;  #10 
a = 8'd50; b = 8'd248;  #10 
a = 8'd50; b = 8'd249;  #10 
a = 8'd50; b = 8'd250;  #10 
a = 8'd50; b = 8'd251;  #10 
a = 8'd50; b = 8'd252;  #10 
a = 8'd50; b = 8'd253;  #10 
a = 8'd50; b = 8'd254;  #10 
a = 8'd50; b = 8'd255;  #10 
a = 8'd51; b = 8'd0;  #10 
a = 8'd51; b = 8'd1;  #10 
a = 8'd51; b = 8'd2;  #10 
a = 8'd51; b = 8'd3;  #10 
a = 8'd51; b = 8'd4;  #10 
a = 8'd51; b = 8'd5;  #10 
a = 8'd51; b = 8'd6;  #10 
a = 8'd51; b = 8'd7;  #10 
a = 8'd51; b = 8'd8;  #10 
a = 8'd51; b = 8'd9;  #10 
a = 8'd51; b = 8'd10;  #10 
a = 8'd51; b = 8'd11;  #10 
a = 8'd51; b = 8'd12;  #10 
a = 8'd51; b = 8'd13;  #10 
a = 8'd51; b = 8'd14;  #10 
a = 8'd51; b = 8'd15;  #10 
a = 8'd51; b = 8'd16;  #10 
a = 8'd51; b = 8'd17;  #10 
a = 8'd51; b = 8'd18;  #10 
a = 8'd51; b = 8'd19;  #10 
a = 8'd51; b = 8'd20;  #10 
a = 8'd51; b = 8'd21;  #10 
a = 8'd51; b = 8'd22;  #10 
a = 8'd51; b = 8'd23;  #10 
a = 8'd51; b = 8'd24;  #10 
a = 8'd51; b = 8'd25;  #10 
a = 8'd51; b = 8'd26;  #10 
a = 8'd51; b = 8'd27;  #10 
a = 8'd51; b = 8'd28;  #10 
a = 8'd51; b = 8'd29;  #10 
a = 8'd51; b = 8'd30;  #10 
a = 8'd51; b = 8'd31;  #10 
a = 8'd51; b = 8'd32;  #10 
a = 8'd51; b = 8'd33;  #10 
a = 8'd51; b = 8'd34;  #10 
a = 8'd51; b = 8'd35;  #10 
a = 8'd51; b = 8'd36;  #10 
a = 8'd51; b = 8'd37;  #10 
a = 8'd51; b = 8'd38;  #10 
a = 8'd51; b = 8'd39;  #10 
a = 8'd51; b = 8'd40;  #10 
a = 8'd51; b = 8'd41;  #10 
a = 8'd51; b = 8'd42;  #10 
a = 8'd51; b = 8'd43;  #10 
a = 8'd51; b = 8'd44;  #10 
a = 8'd51; b = 8'd45;  #10 
a = 8'd51; b = 8'd46;  #10 
a = 8'd51; b = 8'd47;  #10 
a = 8'd51; b = 8'd48;  #10 
a = 8'd51; b = 8'd49;  #10 
a = 8'd51; b = 8'd50;  #10 
a = 8'd51; b = 8'd51;  #10 
a = 8'd51; b = 8'd52;  #10 
a = 8'd51; b = 8'd53;  #10 
a = 8'd51; b = 8'd54;  #10 
a = 8'd51; b = 8'd55;  #10 
a = 8'd51; b = 8'd56;  #10 
a = 8'd51; b = 8'd57;  #10 
a = 8'd51; b = 8'd58;  #10 
a = 8'd51; b = 8'd59;  #10 
a = 8'd51; b = 8'd60;  #10 
a = 8'd51; b = 8'd61;  #10 
a = 8'd51; b = 8'd62;  #10 
a = 8'd51; b = 8'd63;  #10 
a = 8'd51; b = 8'd64;  #10 
a = 8'd51; b = 8'd65;  #10 
a = 8'd51; b = 8'd66;  #10 
a = 8'd51; b = 8'd67;  #10 
a = 8'd51; b = 8'd68;  #10 
a = 8'd51; b = 8'd69;  #10 
a = 8'd51; b = 8'd70;  #10 
a = 8'd51; b = 8'd71;  #10 
a = 8'd51; b = 8'd72;  #10 
a = 8'd51; b = 8'd73;  #10 
a = 8'd51; b = 8'd74;  #10 
a = 8'd51; b = 8'd75;  #10 
a = 8'd51; b = 8'd76;  #10 
a = 8'd51; b = 8'd77;  #10 
a = 8'd51; b = 8'd78;  #10 
a = 8'd51; b = 8'd79;  #10 
a = 8'd51; b = 8'd80;  #10 
a = 8'd51; b = 8'd81;  #10 
a = 8'd51; b = 8'd82;  #10 
a = 8'd51; b = 8'd83;  #10 
a = 8'd51; b = 8'd84;  #10 
a = 8'd51; b = 8'd85;  #10 
a = 8'd51; b = 8'd86;  #10 
a = 8'd51; b = 8'd87;  #10 
a = 8'd51; b = 8'd88;  #10 
a = 8'd51; b = 8'd89;  #10 
a = 8'd51; b = 8'd90;  #10 
a = 8'd51; b = 8'd91;  #10 
a = 8'd51; b = 8'd92;  #10 
a = 8'd51; b = 8'd93;  #10 
a = 8'd51; b = 8'd94;  #10 
a = 8'd51; b = 8'd95;  #10 
a = 8'd51; b = 8'd96;  #10 
a = 8'd51; b = 8'd97;  #10 
a = 8'd51; b = 8'd98;  #10 
a = 8'd51; b = 8'd99;  #10 
a = 8'd51; b = 8'd100;  #10 
a = 8'd51; b = 8'd101;  #10 
a = 8'd51; b = 8'd102;  #10 
a = 8'd51; b = 8'd103;  #10 
a = 8'd51; b = 8'd104;  #10 
a = 8'd51; b = 8'd105;  #10 
a = 8'd51; b = 8'd106;  #10 
a = 8'd51; b = 8'd107;  #10 
a = 8'd51; b = 8'd108;  #10 
a = 8'd51; b = 8'd109;  #10 
a = 8'd51; b = 8'd110;  #10 
a = 8'd51; b = 8'd111;  #10 
a = 8'd51; b = 8'd112;  #10 
a = 8'd51; b = 8'd113;  #10 
a = 8'd51; b = 8'd114;  #10 
a = 8'd51; b = 8'd115;  #10 
a = 8'd51; b = 8'd116;  #10 
a = 8'd51; b = 8'd117;  #10 
a = 8'd51; b = 8'd118;  #10 
a = 8'd51; b = 8'd119;  #10 
a = 8'd51; b = 8'd120;  #10 
a = 8'd51; b = 8'd121;  #10 
a = 8'd51; b = 8'd122;  #10 
a = 8'd51; b = 8'd123;  #10 
a = 8'd51; b = 8'd124;  #10 
a = 8'd51; b = 8'd125;  #10 
a = 8'd51; b = 8'd126;  #10 
a = 8'd51; b = 8'd127;  #10 
a = 8'd51; b = 8'd128;  #10 
a = 8'd51; b = 8'd129;  #10 
a = 8'd51; b = 8'd130;  #10 
a = 8'd51; b = 8'd131;  #10 
a = 8'd51; b = 8'd132;  #10 
a = 8'd51; b = 8'd133;  #10 
a = 8'd51; b = 8'd134;  #10 
a = 8'd51; b = 8'd135;  #10 
a = 8'd51; b = 8'd136;  #10 
a = 8'd51; b = 8'd137;  #10 
a = 8'd51; b = 8'd138;  #10 
a = 8'd51; b = 8'd139;  #10 
a = 8'd51; b = 8'd140;  #10 
a = 8'd51; b = 8'd141;  #10 
a = 8'd51; b = 8'd142;  #10 
a = 8'd51; b = 8'd143;  #10 
a = 8'd51; b = 8'd144;  #10 
a = 8'd51; b = 8'd145;  #10 
a = 8'd51; b = 8'd146;  #10 
a = 8'd51; b = 8'd147;  #10 
a = 8'd51; b = 8'd148;  #10 
a = 8'd51; b = 8'd149;  #10 
a = 8'd51; b = 8'd150;  #10 
a = 8'd51; b = 8'd151;  #10 
a = 8'd51; b = 8'd152;  #10 
a = 8'd51; b = 8'd153;  #10 
a = 8'd51; b = 8'd154;  #10 
a = 8'd51; b = 8'd155;  #10 
a = 8'd51; b = 8'd156;  #10 
a = 8'd51; b = 8'd157;  #10 
a = 8'd51; b = 8'd158;  #10 
a = 8'd51; b = 8'd159;  #10 
a = 8'd51; b = 8'd160;  #10 
a = 8'd51; b = 8'd161;  #10 
a = 8'd51; b = 8'd162;  #10 
a = 8'd51; b = 8'd163;  #10 
a = 8'd51; b = 8'd164;  #10 
a = 8'd51; b = 8'd165;  #10 
a = 8'd51; b = 8'd166;  #10 
a = 8'd51; b = 8'd167;  #10 
a = 8'd51; b = 8'd168;  #10 
a = 8'd51; b = 8'd169;  #10 
a = 8'd51; b = 8'd170;  #10 
a = 8'd51; b = 8'd171;  #10 
a = 8'd51; b = 8'd172;  #10 
a = 8'd51; b = 8'd173;  #10 
a = 8'd51; b = 8'd174;  #10 
a = 8'd51; b = 8'd175;  #10 
a = 8'd51; b = 8'd176;  #10 
a = 8'd51; b = 8'd177;  #10 
a = 8'd51; b = 8'd178;  #10 
a = 8'd51; b = 8'd179;  #10 
a = 8'd51; b = 8'd180;  #10 
a = 8'd51; b = 8'd181;  #10 
a = 8'd51; b = 8'd182;  #10 
a = 8'd51; b = 8'd183;  #10 
a = 8'd51; b = 8'd184;  #10 
a = 8'd51; b = 8'd185;  #10 
a = 8'd51; b = 8'd186;  #10 
a = 8'd51; b = 8'd187;  #10 
a = 8'd51; b = 8'd188;  #10 
a = 8'd51; b = 8'd189;  #10 
a = 8'd51; b = 8'd190;  #10 
a = 8'd51; b = 8'd191;  #10 
a = 8'd51; b = 8'd192;  #10 
a = 8'd51; b = 8'd193;  #10 
a = 8'd51; b = 8'd194;  #10 
a = 8'd51; b = 8'd195;  #10 
a = 8'd51; b = 8'd196;  #10 
a = 8'd51; b = 8'd197;  #10 
a = 8'd51; b = 8'd198;  #10 
a = 8'd51; b = 8'd199;  #10 
a = 8'd51; b = 8'd200;  #10 
a = 8'd51; b = 8'd201;  #10 
a = 8'd51; b = 8'd202;  #10 
a = 8'd51; b = 8'd203;  #10 
a = 8'd51; b = 8'd204;  #10 
a = 8'd51; b = 8'd205;  #10 
a = 8'd51; b = 8'd206;  #10 
a = 8'd51; b = 8'd207;  #10 
a = 8'd51; b = 8'd208;  #10 
a = 8'd51; b = 8'd209;  #10 
a = 8'd51; b = 8'd210;  #10 
a = 8'd51; b = 8'd211;  #10 
a = 8'd51; b = 8'd212;  #10 
a = 8'd51; b = 8'd213;  #10 
a = 8'd51; b = 8'd214;  #10 
a = 8'd51; b = 8'd215;  #10 
a = 8'd51; b = 8'd216;  #10 
a = 8'd51; b = 8'd217;  #10 
a = 8'd51; b = 8'd218;  #10 
a = 8'd51; b = 8'd219;  #10 
a = 8'd51; b = 8'd220;  #10 
a = 8'd51; b = 8'd221;  #10 
a = 8'd51; b = 8'd222;  #10 
a = 8'd51; b = 8'd223;  #10 
a = 8'd51; b = 8'd224;  #10 
a = 8'd51; b = 8'd225;  #10 
a = 8'd51; b = 8'd226;  #10 
a = 8'd51; b = 8'd227;  #10 
a = 8'd51; b = 8'd228;  #10 
a = 8'd51; b = 8'd229;  #10 
a = 8'd51; b = 8'd230;  #10 
a = 8'd51; b = 8'd231;  #10 
a = 8'd51; b = 8'd232;  #10 
a = 8'd51; b = 8'd233;  #10 
a = 8'd51; b = 8'd234;  #10 
a = 8'd51; b = 8'd235;  #10 
a = 8'd51; b = 8'd236;  #10 
a = 8'd51; b = 8'd237;  #10 
a = 8'd51; b = 8'd238;  #10 
a = 8'd51; b = 8'd239;  #10 
a = 8'd51; b = 8'd240;  #10 
a = 8'd51; b = 8'd241;  #10 
a = 8'd51; b = 8'd242;  #10 
a = 8'd51; b = 8'd243;  #10 
a = 8'd51; b = 8'd244;  #10 
a = 8'd51; b = 8'd245;  #10 
a = 8'd51; b = 8'd246;  #10 
a = 8'd51; b = 8'd247;  #10 
a = 8'd51; b = 8'd248;  #10 
a = 8'd51; b = 8'd249;  #10 
a = 8'd51; b = 8'd250;  #10 
a = 8'd51; b = 8'd251;  #10 
a = 8'd51; b = 8'd252;  #10 
a = 8'd51; b = 8'd253;  #10 
a = 8'd51; b = 8'd254;  #10 
a = 8'd51; b = 8'd255;  #10 
a = 8'd52; b = 8'd0;  #10 
a = 8'd52; b = 8'd1;  #10 
a = 8'd52; b = 8'd2;  #10 
a = 8'd52; b = 8'd3;  #10 
a = 8'd52; b = 8'd4;  #10 
a = 8'd52; b = 8'd5;  #10 
a = 8'd52; b = 8'd6;  #10 
a = 8'd52; b = 8'd7;  #10 
a = 8'd52; b = 8'd8;  #10 
a = 8'd52; b = 8'd9;  #10 
a = 8'd52; b = 8'd10;  #10 
a = 8'd52; b = 8'd11;  #10 
a = 8'd52; b = 8'd12;  #10 
a = 8'd52; b = 8'd13;  #10 
a = 8'd52; b = 8'd14;  #10 
a = 8'd52; b = 8'd15;  #10 
a = 8'd52; b = 8'd16;  #10 
a = 8'd52; b = 8'd17;  #10 
a = 8'd52; b = 8'd18;  #10 
a = 8'd52; b = 8'd19;  #10 
a = 8'd52; b = 8'd20;  #10 
a = 8'd52; b = 8'd21;  #10 
a = 8'd52; b = 8'd22;  #10 
a = 8'd52; b = 8'd23;  #10 
a = 8'd52; b = 8'd24;  #10 
a = 8'd52; b = 8'd25;  #10 
a = 8'd52; b = 8'd26;  #10 
a = 8'd52; b = 8'd27;  #10 
a = 8'd52; b = 8'd28;  #10 
a = 8'd52; b = 8'd29;  #10 
a = 8'd52; b = 8'd30;  #10 
a = 8'd52; b = 8'd31;  #10 
a = 8'd52; b = 8'd32;  #10 
a = 8'd52; b = 8'd33;  #10 
a = 8'd52; b = 8'd34;  #10 
a = 8'd52; b = 8'd35;  #10 
a = 8'd52; b = 8'd36;  #10 
a = 8'd52; b = 8'd37;  #10 
a = 8'd52; b = 8'd38;  #10 
a = 8'd52; b = 8'd39;  #10 
a = 8'd52; b = 8'd40;  #10 
a = 8'd52; b = 8'd41;  #10 
a = 8'd52; b = 8'd42;  #10 
a = 8'd52; b = 8'd43;  #10 
a = 8'd52; b = 8'd44;  #10 
a = 8'd52; b = 8'd45;  #10 
a = 8'd52; b = 8'd46;  #10 
a = 8'd52; b = 8'd47;  #10 
a = 8'd52; b = 8'd48;  #10 
a = 8'd52; b = 8'd49;  #10 
a = 8'd52; b = 8'd50;  #10 
a = 8'd52; b = 8'd51;  #10 
a = 8'd52; b = 8'd52;  #10 
a = 8'd52; b = 8'd53;  #10 
a = 8'd52; b = 8'd54;  #10 
a = 8'd52; b = 8'd55;  #10 
a = 8'd52; b = 8'd56;  #10 
a = 8'd52; b = 8'd57;  #10 
a = 8'd52; b = 8'd58;  #10 
a = 8'd52; b = 8'd59;  #10 
a = 8'd52; b = 8'd60;  #10 
a = 8'd52; b = 8'd61;  #10 
a = 8'd52; b = 8'd62;  #10 
a = 8'd52; b = 8'd63;  #10 
a = 8'd52; b = 8'd64;  #10 
a = 8'd52; b = 8'd65;  #10 
a = 8'd52; b = 8'd66;  #10 
a = 8'd52; b = 8'd67;  #10 
a = 8'd52; b = 8'd68;  #10 
a = 8'd52; b = 8'd69;  #10 
a = 8'd52; b = 8'd70;  #10 
a = 8'd52; b = 8'd71;  #10 
a = 8'd52; b = 8'd72;  #10 
a = 8'd52; b = 8'd73;  #10 
a = 8'd52; b = 8'd74;  #10 
a = 8'd52; b = 8'd75;  #10 
a = 8'd52; b = 8'd76;  #10 
a = 8'd52; b = 8'd77;  #10 
a = 8'd52; b = 8'd78;  #10 
a = 8'd52; b = 8'd79;  #10 
a = 8'd52; b = 8'd80;  #10 
a = 8'd52; b = 8'd81;  #10 
a = 8'd52; b = 8'd82;  #10 
a = 8'd52; b = 8'd83;  #10 
a = 8'd52; b = 8'd84;  #10 
a = 8'd52; b = 8'd85;  #10 
a = 8'd52; b = 8'd86;  #10 
a = 8'd52; b = 8'd87;  #10 
a = 8'd52; b = 8'd88;  #10 
a = 8'd52; b = 8'd89;  #10 
a = 8'd52; b = 8'd90;  #10 
a = 8'd52; b = 8'd91;  #10 
a = 8'd52; b = 8'd92;  #10 
a = 8'd52; b = 8'd93;  #10 
a = 8'd52; b = 8'd94;  #10 
a = 8'd52; b = 8'd95;  #10 
a = 8'd52; b = 8'd96;  #10 
a = 8'd52; b = 8'd97;  #10 
a = 8'd52; b = 8'd98;  #10 
a = 8'd52; b = 8'd99;  #10 
a = 8'd52; b = 8'd100;  #10 
a = 8'd52; b = 8'd101;  #10 
a = 8'd52; b = 8'd102;  #10 
a = 8'd52; b = 8'd103;  #10 
a = 8'd52; b = 8'd104;  #10 
a = 8'd52; b = 8'd105;  #10 
a = 8'd52; b = 8'd106;  #10 
a = 8'd52; b = 8'd107;  #10 
a = 8'd52; b = 8'd108;  #10 
a = 8'd52; b = 8'd109;  #10 
a = 8'd52; b = 8'd110;  #10 
a = 8'd52; b = 8'd111;  #10 
a = 8'd52; b = 8'd112;  #10 
a = 8'd52; b = 8'd113;  #10 
a = 8'd52; b = 8'd114;  #10 
a = 8'd52; b = 8'd115;  #10 
a = 8'd52; b = 8'd116;  #10 
a = 8'd52; b = 8'd117;  #10 
a = 8'd52; b = 8'd118;  #10 
a = 8'd52; b = 8'd119;  #10 
a = 8'd52; b = 8'd120;  #10 
a = 8'd52; b = 8'd121;  #10 
a = 8'd52; b = 8'd122;  #10 
a = 8'd52; b = 8'd123;  #10 
a = 8'd52; b = 8'd124;  #10 
a = 8'd52; b = 8'd125;  #10 
a = 8'd52; b = 8'd126;  #10 
a = 8'd52; b = 8'd127;  #10 
a = 8'd52; b = 8'd128;  #10 
a = 8'd52; b = 8'd129;  #10 
a = 8'd52; b = 8'd130;  #10 
a = 8'd52; b = 8'd131;  #10 
a = 8'd52; b = 8'd132;  #10 
a = 8'd52; b = 8'd133;  #10 
a = 8'd52; b = 8'd134;  #10 
a = 8'd52; b = 8'd135;  #10 
a = 8'd52; b = 8'd136;  #10 
a = 8'd52; b = 8'd137;  #10 
a = 8'd52; b = 8'd138;  #10 
a = 8'd52; b = 8'd139;  #10 
a = 8'd52; b = 8'd140;  #10 
a = 8'd52; b = 8'd141;  #10 
a = 8'd52; b = 8'd142;  #10 
a = 8'd52; b = 8'd143;  #10 
a = 8'd52; b = 8'd144;  #10 
a = 8'd52; b = 8'd145;  #10 
a = 8'd52; b = 8'd146;  #10 
a = 8'd52; b = 8'd147;  #10 
a = 8'd52; b = 8'd148;  #10 
a = 8'd52; b = 8'd149;  #10 
a = 8'd52; b = 8'd150;  #10 
a = 8'd52; b = 8'd151;  #10 
a = 8'd52; b = 8'd152;  #10 
a = 8'd52; b = 8'd153;  #10 
a = 8'd52; b = 8'd154;  #10 
a = 8'd52; b = 8'd155;  #10 
a = 8'd52; b = 8'd156;  #10 
a = 8'd52; b = 8'd157;  #10 
a = 8'd52; b = 8'd158;  #10 
a = 8'd52; b = 8'd159;  #10 
a = 8'd52; b = 8'd160;  #10 
a = 8'd52; b = 8'd161;  #10 
a = 8'd52; b = 8'd162;  #10 
a = 8'd52; b = 8'd163;  #10 
a = 8'd52; b = 8'd164;  #10 
a = 8'd52; b = 8'd165;  #10 
a = 8'd52; b = 8'd166;  #10 
a = 8'd52; b = 8'd167;  #10 
a = 8'd52; b = 8'd168;  #10 
a = 8'd52; b = 8'd169;  #10 
a = 8'd52; b = 8'd170;  #10 
a = 8'd52; b = 8'd171;  #10 
a = 8'd52; b = 8'd172;  #10 
a = 8'd52; b = 8'd173;  #10 
a = 8'd52; b = 8'd174;  #10 
a = 8'd52; b = 8'd175;  #10 
a = 8'd52; b = 8'd176;  #10 
a = 8'd52; b = 8'd177;  #10 
a = 8'd52; b = 8'd178;  #10 
a = 8'd52; b = 8'd179;  #10 
a = 8'd52; b = 8'd180;  #10 
a = 8'd52; b = 8'd181;  #10 
a = 8'd52; b = 8'd182;  #10 
a = 8'd52; b = 8'd183;  #10 
a = 8'd52; b = 8'd184;  #10 
a = 8'd52; b = 8'd185;  #10 
a = 8'd52; b = 8'd186;  #10 
a = 8'd52; b = 8'd187;  #10 
a = 8'd52; b = 8'd188;  #10 
a = 8'd52; b = 8'd189;  #10 
a = 8'd52; b = 8'd190;  #10 
a = 8'd52; b = 8'd191;  #10 
a = 8'd52; b = 8'd192;  #10 
a = 8'd52; b = 8'd193;  #10 
a = 8'd52; b = 8'd194;  #10 
a = 8'd52; b = 8'd195;  #10 
a = 8'd52; b = 8'd196;  #10 
a = 8'd52; b = 8'd197;  #10 
a = 8'd52; b = 8'd198;  #10 
a = 8'd52; b = 8'd199;  #10 
a = 8'd52; b = 8'd200;  #10 
a = 8'd52; b = 8'd201;  #10 
a = 8'd52; b = 8'd202;  #10 
a = 8'd52; b = 8'd203;  #10 
a = 8'd52; b = 8'd204;  #10 
a = 8'd52; b = 8'd205;  #10 
a = 8'd52; b = 8'd206;  #10 
a = 8'd52; b = 8'd207;  #10 
a = 8'd52; b = 8'd208;  #10 
a = 8'd52; b = 8'd209;  #10 
a = 8'd52; b = 8'd210;  #10 
a = 8'd52; b = 8'd211;  #10 
a = 8'd52; b = 8'd212;  #10 
a = 8'd52; b = 8'd213;  #10 
a = 8'd52; b = 8'd214;  #10 
a = 8'd52; b = 8'd215;  #10 
a = 8'd52; b = 8'd216;  #10 
a = 8'd52; b = 8'd217;  #10 
a = 8'd52; b = 8'd218;  #10 
a = 8'd52; b = 8'd219;  #10 
a = 8'd52; b = 8'd220;  #10 
a = 8'd52; b = 8'd221;  #10 
a = 8'd52; b = 8'd222;  #10 
a = 8'd52; b = 8'd223;  #10 
a = 8'd52; b = 8'd224;  #10 
a = 8'd52; b = 8'd225;  #10 
a = 8'd52; b = 8'd226;  #10 
a = 8'd52; b = 8'd227;  #10 
a = 8'd52; b = 8'd228;  #10 
a = 8'd52; b = 8'd229;  #10 
a = 8'd52; b = 8'd230;  #10 
a = 8'd52; b = 8'd231;  #10 
a = 8'd52; b = 8'd232;  #10 
a = 8'd52; b = 8'd233;  #10 
a = 8'd52; b = 8'd234;  #10 
a = 8'd52; b = 8'd235;  #10 
a = 8'd52; b = 8'd236;  #10 
a = 8'd52; b = 8'd237;  #10 
a = 8'd52; b = 8'd238;  #10 
a = 8'd52; b = 8'd239;  #10 
a = 8'd52; b = 8'd240;  #10 
a = 8'd52; b = 8'd241;  #10 
a = 8'd52; b = 8'd242;  #10 
a = 8'd52; b = 8'd243;  #10 
a = 8'd52; b = 8'd244;  #10 
a = 8'd52; b = 8'd245;  #10 
a = 8'd52; b = 8'd246;  #10 
a = 8'd52; b = 8'd247;  #10 
a = 8'd52; b = 8'd248;  #10 
a = 8'd52; b = 8'd249;  #10 
a = 8'd52; b = 8'd250;  #10 
a = 8'd52; b = 8'd251;  #10 
a = 8'd52; b = 8'd252;  #10 
a = 8'd52; b = 8'd253;  #10 
a = 8'd52; b = 8'd254;  #10 
a = 8'd52; b = 8'd255;  #10 
a = 8'd53; b = 8'd0;  #10 
a = 8'd53; b = 8'd1;  #10 
a = 8'd53; b = 8'd2;  #10 
a = 8'd53; b = 8'd3;  #10 
a = 8'd53; b = 8'd4;  #10 
a = 8'd53; b = 8'd5;  #10 
a = 8'd53; b = 8'd6;  #10 
a = 8'd53; b = 8'd7;  #10 
a = 8'd53; b = 8'd8;  #10 
a = 8'd53; b = 8'd9;  #10 
a = 8'd53; b = 8'd10;  #10 
a = 8'd53; b = 8'd11;  #10 
a = 8'd53; b = 8'd12;  #10 
a = 8'd53; b = 8'd13;  #10 
a = 8'd53; b = 8'd14;  #10 
a = 8'd53; b = 8'd15;  #10 
a = 8'd53; b = 8'd16;  #10 
a = 8'd53; b = 8'd17;  #10 
a = 8'd53; b = 8'd18;  #10 
a = 8'd53; b = 8'd19;  #10 
a = 8'd53; b = 8'd20;  #10 
a = 8'd53; b = 8'd21;  #10 
a = 8'd53; b = 8'd22;  #10 
a = 8'd53; b = 8'd23;  #10 
a = 8'd53; b = 8'd24;  #10 
a = 8'd53; b = 8'd25;  #10 
a = 8'd53; b = 8'd26;  #10 
a = 8'd53; b = 8'd27;  #10 
a = 8'd53; b = 8'd28;  #10 
a = 8'd53; b = 8'd29;  #10 
a = 8'd53; b = 8'd30;  #10 
a = 8'd53; b = 8'd31;  #10 
a = 8'd53; b = 8'd32;  #10 
a = 8'd53; b = 8'd33;  #10 
a = 8'd53; b = 8'd34;  #10 
a = 8'd53; b = 8'd35;  #10 
a = 8'd53; b = 8'd36;  #10 
a = 8'd53; b = 8'd37;  #10 
a = 8'd53; b = 8'd38;  #10 
a = 8'd53; b = 8'd39;  #10 
a = 8'd53; b = 8'd40;  #10 
a = 8'd53; b = 8'd41;  #10 
a = 8'd53; b = 8'd42;  #10 
a = 8'd53; b = 8'd43;  #10 
a = 8'd53; b = 8'd44;  #10 
a = 8'd53; b = 8'd45;  #10 
a = 8'd53; b = 8'd46;  #10 
a = 8'd53; b = 8'd47;  #10 
a = 8'd53; b = 8'd48;  #10 
a = 8'd53; b = 8'd49;  #10 
a = 8'd53; b = 8'd50;  #10 
a = 8'd53; b = 8'd51;  #10 
a = 8'd53; b = 8'd52;  #10 
a = 8'd53; b = 8'd53;  #10 
a = 8'd53; b = 8'd54;  #10 
a = 8'd53; b = 8'd55;  #10 
a = 8'd53; b = 8'd56;  #10 
a = 8'd53; b = 8'd57;  #10 
a = 8'd53; b = 8'd58;  #10 
a = 8'd53; b = 8'd59;  #10 
a = 8'd53; b = 8'd60;  #10 
a = 8'd53; b = 8'd61;  #10 
a = 8'd53; b = 8'd62;  #10 
a = 8'd53; b = 8'd63;  #10 
a = 8'd53; b = 8'd64;  #10 
a = 8'd53; b = 8'd65;  #10 
a = 8'd53; b = 8'd66;  #10 
a = 8'd53; b = 8'd67;  #10 
a = 8'd53; b = 8'd68;  #10 
a = 8'd53; b = 8'd69;  #10 
a = 8'd53; b = 8'd70;  #10 
a = 8'd53; b = 8'd71;  #10 
a = 8'd53; b = 8'd72;  #10 
a = 8'd53; b = 8'd73;  #10 
a = 8'd53; b = 8'd74;  #10 
a = 8'd53; b = 8'd75;  #10 
a = 8'd53; b = 8'd76;  #10 
a = 8'd53; b = 8'd77;  #10 
a = 8'd53; b = 8'd78;  #10 
a = 8'd53; b = 8'd79;  #10 
a = 8'd53; b = 8'd80;  #10 
a = 8'd53; b = 8'd81;  #10 
a = 8'd53; b = 8'd82;  #10 
a = 8'd53; b = 8'd83;  #10 
a = 8'd53; b = 8'd84;  #10 
a = 8'd53; b = 8'd85;  #10 
a = 8'd53; b = 8'd86;  #10 
a = 8'd53; b = 8'd87;  #10 
a = 8'd53; b = 8'd88;  #10 
a = 8'd53; b = 8'd89;  #10 
a = 8'd53; b = 8'd90;  #10 
a = 8'd53; b = 8'd91;  #10 
a = 8'd53; b = 8'd92;  #10 
a = 8'd53; b = 8'd93;  #10 
a = 8'd53; b = 8'd94;  #10 
a = 8'd53; b = 8'd95;  #10 
a = 8'd53; b = 8'd96;  #10 
a = 8'd53; b = 8'd97;  #10 
a = 8'd53; b = 8'd98;  #10 
a = 8'd53; b = 8'd99;  #10 
a = 8'd53; b = 8'd100;  #10 
a = 8'd53; b = 8'd101;  #10 
a = 8'd53; b = 8'd102;  #10 
a = 8'd53; b = 8'd103;  #10 
a = 8'd53; b = 8'd104;  #10 
a = 8'd53; b = 8'd105;  #10 
a = 8'd53; b = 8'd106;  #10 
a = 8'd53; b = 8'd107;  #10 
a = 8'd53; b = 8'd108;  #10 
a = 8'd53; b = 8'd109;  #10 
a = 8'd53; b = 8'd110;  #10 
a = 8'd53; b = 8'd111;  #10 
a = 8'd53; b = 8'd112;  #10 
a = 8'd53; b = 8'd113;  #10 
a = 8'd53; b = 8'd114;  #10 
a = 8'd53; b = 8'd115;  #10 
a = 8'd53; b = 8'd116;  #10 
a = 8'd53; b = 8'd117;  #10 
a = 8'd53; b = 8'd118;  #10 
a = 8'd53; b = 8'd119;  #10 
a = 8'd53; b = 8'd120;  #10 
a = 8'd53; b = 8'd121;  #10 
a = 8'd53; b = 8'd122;  #10 
a = 8'd53; b = 8'd123;  #10 
a = 8'd53; b = 8'd124;  #10 
a = 8'd53; b = 8'd125;  #10 
a = 8'd53; b = 8'd126;  #10 
a = 8'd53; b = 8'd127;  #10 
a = 8'd53; b = 8'd128;  #10 
a = 8'd53; b = 8'd129;  #10 
a = 8'd53; b = 8'd130;  #10 
a = 8'd53; b = 8'd131;  #10 
a = 8'd53; b = 8'd132;  #10 
a = 8'd53; b = 8'd133;  #10 
a = 8'd53; b = 8'd134;  #10 
a = 8'd53; b = 8'd135;  #10 
a = 8'd53; b = 8'd136;  #10 
a = 8'd53; b = 8'd137;  #10 
a = 8'd53; b = 8'd138;  #10 
a = 8'd53; b = 8'd139;  #10 
a = 8'd53; b = 8'd140;  #10 
a = 8'd53; b = 8'd141;  #10 
a = 8'd53; b = 8'd142;  #10 
a = 8'd53; b = 8'd143;  #10 
a = 8'd53; b = 8'd144;  #10 
a = 8'd53; b = 8'd145;  #10 
a = 8'd53; b = 8'd146;  #10 
a = 8'd53; b = 8'd147;  #10 
a = 8'd53; b = 8'd148;  #10 
a = 8'd53; b = 8'd149;  #10 
a = 8'd53; b = 8'd150;  #10 
a = 8'd53; b = 8'd151;  #10 
a = 8'd53; b = 8'd152;  #10 
a = 8'd53; b = 8'd153;  #10 
a = 8'd53; b = 8'd154;  #10 
a = 8'd53; b = 8'd155;  #10 
a = 8'd53; b = 8'd156;  #10 
a = 8'd53; b = 8'd157;  #10 
a = 8'd53; b = 8'd158;  #10 
a = 8'd53; b = 8'd159;  #10 
a = 8'd53; b = 8'd160;  #10 
a = 8'd53; b = 8'd161;  #10 
a = 8'd53; b = 8'd162;  #10 
a = 8'd53; b = 8'd163;  #10 
a = 8'd53; b = 8'd164;  #10 
a = 8'd53; b = 8'd165;  #10 
a = 8'd53; b = 8'd166;  #10 
a = 8'd53; b = 8'd167;  #10 
a = 8'd53; b = 8'd168;  #10 
a = 8'd53; b = 8'd169;  #10 
a = 8'd53; b = 8'd170;  #10 
a = 8'd53; b = 8'd171;  #10 
a = 8'd53; b = 8'd172;  #10 
a = 8'd53; b = 8'd173;  #10 
a = 8'd53; b = 8'd174;  #10 
a = 8'd53; b = 8'd175;  #10 
a = 8'd53; b = 8'd176;  #10 
a = 8'd53; b = 8'd177;  #10 
a = 8'd53; b = 8'd178;  #10 
a = 8'd53; b = 8'd179;  #10 
a = 8'd53; b = 8'd180;  #10 
a = 8'd53; b = 8'd181;  #10 
a = 8'd53; b = 8'd182;  #10 
a = 8'd53; b = 8'd183;  #10 
a = 8'd53; b = 8'd184;  #10 
a = 8'd53; b = 8'd185;  #10 
a = 8'd53; b = 8'd186;  #10 
a = 8'd53; b = 8'd187;  #10 
a = 8'd53; b = 8'd188;  #10 
a = 8'd53; b = 8'd189;  #10 
a = 8'd53; b = 8'd190;  #10 
a = 8'd53; b = 8'd191;  #10 
a = 8'd53; b = 8'd192;  #10 
a = 8'd53; b = 8'd193;  #10 
a = 8'd53; b = 8'd194;  #10 
a = 8'd53; b = 8'd195;  #10 
a = 8'd53; b = 8'd196;  #10 
a = 8'd53; b = 8'd197;  #10 
a = 8'd53; b = 8'd198;  #10 
a = 8'd53; b = 8'd199;  #10 
a = 8'd53; b = 8'd200;  #10 
a = 8'd53; b = 8'd201;  #10 
a = 8'd53; b = 8'd202;  #10 
a = 8'd53; b = 8'd203;  #10 
a = 8'd53; b = 8'd204;  #10 
a = 8'd53; b = 8'd205;  #10 
a = 8'd53; b = 8'd206;  #10 
a = 8'd53; b = 8'd207;  #10 
a = 8'd53; b = 8'd208;  #10 
a = 8'd53; b = 8'd209;  #10 
a = 8'd53; b = 8'd210;  #10 
a = 8'd53; b = 8'd211;  #10 
a = 8'd53; b = 8'd212;  #10 
a = 8'd53; b = 8'd213;  #10 
a = 8'd53; b = 8'd214;  #10 
a = 8'd53; b = 8'd215;  #10 
a = 8'd53; b = 8'd216;  #10 
a = 8'd53; b = 8'd217;  #10 
a = 8'd53; b = 8'd218;  #10 
a = 8'd53; b = 8'd219;  #10 
a = 8'd53; b = 8'd220;  #10 
a = 8'd53; b = 8'd221;  #10 
a = 8'd53; b = 8'd222;  #10 
a = 8'd53; b = 8'd223;  #10 
a = 8'd53; b = 8'd224;  #10 
a = 8'd53; b = 8'd225;  #10 
a = 8'd53; b = 8'd226;  #10 
a = 8'd53; b = 8'd227;  #10 
a = 8'd53; b = 8'd228;  #10 
a = 8'd53; b = 8'd229;  #10 
a = 8'd53; b = 8'd230;  #10 
a = 8'd53; b = 8'd231;  #10 
a = 8'd53; b = 8'd232;  #10 
a = 8'd53; b = 8'd233;  #10 
a = 8'd53; b = 8'd234;  #10 
a = 8'd53; b = 8'd235;  #10 
a = 8'd53; b = 8'd236;  #10 
a = 8'd53; b = 8'd237;  #10 
a = 8'd53; b = 8'd238;  #10 
a = 8'd53; b = 8'd239;  #10 
a = 8'd53; b = 8'd240;  #10 
a = 8'd53; b = 8'd241;  #10 
a = 8'd53; b = 8'd242;  #10 
a = 8'd53; b = 8'd243;  #10 
a = 8'd53; b = 8'd244;  #10 
a = 8'd53; b = 8'd245;  #10 
a = 8'd53; b = 8'd246;  #10 
a = 8'd53; b = 8'd247;  #10 
a = 8'd53; b = 8'd248;  #10 
a = 8'd53; b = 8'd249;  #10 
a = 8'd53; b = 8'd250;  #10 
a = 8'd53; b = 8'd251;  #10 
a = 8'd53; b = 8'd252;  #10 
a = 8'd53; b = 8'd253;  #10 
a = 8'd53; b = 8'd254;  #10 
a = 8'd53; b = 8'd255;  #10 
a = 8'd54; b = 8'd0;  #10 
a = 8'd54; b = 8'd1;  #10 
a = 8'd54; b = 8'd2;  #10 
a = 8'd54; b = 8'd3;  #10 
a = 8'd54; b = 8'd4;  #10 
a = 8'd54; b = 8'd5;  #10 
a = 8'd54; b = 8'd6;  #10 
a = 8'd54; b = 8'd7;  #10 
a = 8'd54; b = 8'd8;  #10 
a = 8'd54; b = 8'd9;  #10 
a = 8'd54; b = 8'd10;  #10 
a = 8'd54; b = 8'd11;  #10 
a = 8'd54; b = 8'd12;  #10 
a = 8'd54; b = 8'd13;  #10 
a = 8'd54; b = 8'd14;  #10 
a = 8'd54; b = 8'd15;  #10 
a = 8'd54; b = 8'd16;  #10 
a = 8'd54; b = 8'd17;  #10 
a = 8'd54; b = 8'd18;  #10 
a = 8'd54; b = 8'd19;  #10 
a = 8'd54; b = 8'd20;  #10 
a = 8'd54; b = 8'd21;  #10 
a = 8'd54; b = 8'd22;  #10 
a = 8'd54; b = 8'd23;  #10 
a = 8'd54; b = 8'd24;  #10 
a = 8'd54; b = 8'd25;  #10 
a = 8'd54; b = 8'd26;  #10 
a = 8'd54; b = 8'd27;  #10 
a = 8'd54; b = 8'd28;  #10 
a = 8'd54; b = 8'd29;  #10 
a = 8'd54; b = 8'd30;  #10 
a = 8'd54; b = 8'd31;  #10 
a = 8'd54; b = 8'd32;  #10 
a = 8'd54; b = 8'd33;  #10 
a = 8'd54; b = 8'd34;  #10 
a = 8'd54; b = 8'd35;  #10 
a = 8'd54; b = 8'd36;  #10 
a = 8'd54; b = 8'd37;  #10 
a = 8'd54; b = 8'd38;  #10 
a = 8'd54; b = 8'd39;  #10 
a = 8'd54; b = 8'd40;  #10 
a = 8'd54; b = 8'd41;  #10 
a = 8'd54; b = 8'd42;  #10 
a = 8'd54; b = 8'd43;  #10 
a = 8'd54; b = 8'd44;  #10 
a = 8'd54; b = 8'd45;  #10 
a = 8'd54; b = 8'd46;  #10 
a = 8'd54; b = 8'd47;  #10 
a = 8'd54; b = 8'd48;  #10 
a = 8'd54; b = 8'd49;  #10 
a = 8'd54; b = 8'd50;  #10 
a = 8'd54; b = 8'd51;  #10 
a = 8'd54; b = 8'd52;  #10 
a = 8'd54; b = 8'd53;  #10 
a = 8'd54; b = 8'd54;  #10 
a = 8'd54; b = 8'd55;  #10 
a = 8'd54; b = 8'd56;  #10 
a = 8'd54; b = 8'd57;  #10 
a = 8'd54; b = 8'd58;  #10 
a = 8'd54; b = 8'd59;  #10 
a = 8'd54; b = 8'd60;  #10 
a = 8'd54; b = 8'd61;  #10 
a = 8'd54; b = 8'd62;  #10 
a = 8'd54; b = 8'd63;  #10 
a = 8'd54; b = 8'd64;  #10 
a = 8'd54; b = 8'd65;  #10 
a = 8'd54; b = 8'd66;  #10 
a = 8'd54; b = 8'd67;  #10 
a = 8'd54; b = 8'd68;  #10 
a = 8'd54; b = 8'd69;  #10 
a = 8'd54; b = 8'd70;  #10 
a = 8'd54; b = 8'd71;  #10 
a = 8'd54; b = 8'd72;  #10 
a = 8'd54; b = 8'd73;  #10 
a = 8'd54; b = 8'd74;  #10 
a = 8'd54; b = 8'd75;  #10 
a = 8'd54; b = 8'd76;  #10 
a = 8'd54; b = 8'd77;  #10 
a = 8'd54; b = 8'd78;  #10 
a = 8'd54; b = 8'd79;  #10 
a = 8'd54; b = 8'd80;  #10 
a = 8'd54; b = 8'd81;  #10 
a = 8'd54; b = 8'd82;  #10 
a = 8'd54; b = 8'd83;  #10 
a = 8'd54; b = 8'd84;  #10 
a = 8'd54; b = 8'd85;  #10 
a = 8'd54; b = 8'd86;  #10 
a = 8'd54; b = 8'd87;  #10 
a = 8'd54; b = 8'd88;  #10 
a = 8'd54; b = 8'd89;  #10 
a = 8'd54; b = 8'd90;  #10 
a = 8'd54; b = 8'd91;  #10 
a = 8'd54; b = 8'd92;  #10 
a = 8'd54; b = 8'd93;  #10 
a = 8'd54; b = 8'd94;  #10 
a = 8'd54; b = 8'd95;  #10 
a = 8'd54; b = 8'd96;  #10 
a = 8'd54; b = 8'd97;  #10 
a = 8'd54; b = 8'd98;  #10 
a = 8'd54; b = 8'd99;  #10 
a = 8'd54; b = 8'd100;  #10 
a = 8'd54; b = 8'd101;  #10 
a = 8'd54; b = 8'd102;  #10 
a = 8'd54; b = 8'd103;  #10 
a = 8'd54; b = 8'd104;  #10 
a = 8'd54; b = 8'd105;  #10 
a = 8'd54; b = 8'd106;  #10 
a = 8'd54; b = 8'd107;  #10 
a = 8'd54; b = 8'd108;  #10 
a = 8'd54; b = 8'd109;  #10 
a = 8'd54; b = 8'd110;  #10 
a = 8'd54; b = 8'd111;  #10 
a = 8'd54; b = 8'd112;  #10 
a = 8'd54; b = 8'd113;  #10 
a = 8'd54; b = 8'd114;  #10 
a = 8'd54; b = 8'd115;  #10 
a = 8'd54; b = 8'd116;  #10 
a = 8'd54; b = 8'd117;  #10 
a = 8'd54; b = 8'd118;  #10 
a = 8'd54; b = 8'd119;  #10 
a = 8'd54; b = 8'd120;  #10 
a = 8'd54; b = 8'd121;  #10 
a = 8'd54; b = 8'd122;  #10 
a = 8'd54; b = 8'd123;  #10 
a = 8'd54; b = 8'd124;  #10 
a = 8'd54; b = 8'd125;  #10 
a = 8'd54; b = 8'd126;  #10 
a = 8'd54; b = 8'd127;  #10 
a = 8'd54; b = 8'd128;  #10 
a = 8'd54; b = 8'd129;  #10 
a = 8'd54; b = 8'd130;  #10 
a = 8'd54; b = 8'd131;  #10 
a = 8'd54; b = 8'd132;  #10 
a = 8'd54; b = 8'd133;  #10 
a = 8'd54; b = 8'd134;  #10 
a = 8'd54; b = 8'd135;  #10 
a = 8'd54; b = 8'd136;  #10 
a = 8'd54; b = 8'd137;  #10 
a = 8'd54; b = 8'd138;  #10 
a = 8'd54; b = 8'd139;  #10 
a = 8'd54; b = 8'd140;  #10 
a = 8'd54; b = 8'd141;  #10 
a = 8'd54; b = 8'd142;  #10 
a = 8'd54; b = 8'd143;  #10 
a = 8'd54; b = 8'd144;  #10 
a = 8'd54; b = 8'd145;  #10 
a = 8'd54; b = 8'd146;  #10 
a = 8'd54; b = 8'd147;  #10 
a = 8'd54; b = 8'd148;  #10 
a = 8'd54; b = 8'd149;  #10 
a = 8'd54; b = 8'd150;  #10 
a = 8'd54; b = 8'd151;  #10 
a = 8'd54; b = 8'd152;  #10 
a = 8'd54; b = 8'd153;  #10 
a = 8'd54; b = 8'd154;  #10 
a = 8'd54; b = 8'd155;  #10 
a = 8'd54; b = 8'd156;  #10 
a = 8'd54; b = 8'd157;  #10 
a = 8'd54; b = 8'd158;  #10 
a = 8'd54; b = 8'd159;  #10 
a = 8'd54; b = 8'd160;  #10 
a = 8'd54; b = 8'd161;  #10 
a = 8'd54; b = 8'd162;  #10 
a = 8'd54; b = 8'd163;  #10 
a = 8'd54; b = 8'd164;  #10 
a = 8'd54; b = 8'd165;  #10 
a = 8'd54; b = 8'd166;  #10 
a = 8'd54; b = 8'd167;  #10 
a = 8'd54; b = 8'd168;  #10 
a = 8'd54; b = 8'd169;  #10 
a = 8'd54; b = 8'd170;  #10 
a = 8'd54; b = 8'd171;  #10 
a = 8'd54; b = 8'd172;  #10 
a = 8'd54; b = 8'd173;  #10 
a = 8'd54; b = 8'd174;  #10 
a = 8'd54; b = 8'd175;  #10 
a = 8'd54; b = 8'd176;  #10 
a = 8'd54; b = 8'd177;  #10 
a = 8'd54; b = 8'd178;  #10 
a = 8'd54; b = 8'd179;  #10 
a = 8'd54; b = 8'd180;  #10 
a = 8'd54; b = 8'd181;  #10 
a = 8'd54; b = 8'd182;  #10 
a = 8'd54; b = 8'd183;  #10 
a = 8'd54; b = 8'd184;  #10 
a = 8'd54; b = 8'd185;  #10 
a = 8'd54; b = 8'd186;  #10 
a = 8'd54; b = 8'd187;  #10 
a = 8'd54; b = 8'd188;  #10 
a = 8'd54; b = 8'd189;  #10 
a = 8'd54; b = 8'd190;  #10 
a = 8'd54; b = 8'd191;  #10 
a = 8'd54; b = 8'd192;  #10 
a = 8'd54; b = 8'd193;  #10 
a = 8'd54; b = 8'd194;  #10 
a = 8'd54; b = 8'd195;  #10 
a = 8'd54; b = 8'd196;  #10 
a = 8'd54; b = 8'd197;  #10 
a = 8'd54; b = 8'd198;  #10 
a = 8'd54; b = 8'd199;  #10 
a = 8'd54; b = 8'd200;  #10 
a = 8'd54; b = 8'd201;  #10 
a = 8'd54; b = 8'd202;  #10 
a = 8'd54; b = 8'd203;  #10 
a = 8'd54; b = 8'd204;  #10 
a = 8'd54; b = 8'd205;  #10 
a = 8'd54; b = 8'd206;  #10 
a = 8'd54; b = 8'd207;  #10 
a = 8'd54; b = 8'd208;  #10 
a = 8'd54; b = 8'd209;  #10 
a = 8'd54; b = 8'd210;  #10 
a = 8'd54; b = 8'd211;  #10 
a = 8'd54; b = 8'd212;  #10 
a = 8'd54; b = 8'd213;  #10 
a = 8'd54; b = 8'd214;  #10 
a = 8'd54; b = 8'd215;  #10 
a = 8'd54; b = 8'd216;  #10 
a = 8'd54; b = 8'd217;  #10 
a = 8'd54; b = 8'd218;  #10 
a = 8'd54; b = 8'd219;  #10 
a = 8'd54; b = 8'd220;  #10 
a = 8'd54; b = 8'd221;  #10 
a = 8'd54; b = 8'd222;  #10 
a = 8'd54; b = 8'd223;  #10 
a = 8'd54; b = 8'd224;  #10 
a = 8'd54; b = 8'd225;  #10 
a = 8'd54; b = 8'd226;  #10 
a = 8'd54; b = 8'd227;  #10 
a = 8'd54; b = 8'd228;  #10 
a = 8'd54; b = 8'd229;  #10 
a = 8'd54; b = 8'd230;  #10 
a = 8'd54; b = 8'd231;  #10 
a = 8'd54; b = 8'd232;  #10 
a = 8'd54; b = 8'd233;  #10 
a = 8'd54; b = 8'd234;  #10 
a = 8'd54; b = 8'd235;  #10 
a = 8'd54; b = 8'd236;  #10 
a = 8'd54; b = 8'd237;  #10 
a = 8'd54; b = 8'd238;  #10 
a = 8'd54; b = 8'd239;  #10 
a = 8'd54; b = 8'd240;  #10 
a = 8'd54; b = 8'd241;  #10 
a = 8'd54; b = 8'd242;  #10 
a = 8'd54; b = 8'd243;  #10 
a = 8'd54; b = 8'd244;  #10 
a = 8'd54; b = 8'd245;  #10 
a = 8'd54; b = 8'd246;  #10 
a = 8'd54; b = 8'd247;  #10 
a = 8'd54; b = 8'd248;  #10 
a = 8'd54; b = 8'd249;  #10 
a = 8'd54; b = 8'd250;  #10 
a = 8'd54; b = 8'd251;  #10 
a = 8'd54; b = 8'd252;  #10 
a = 8'd54; b = 8'd253;  #10 
a = 8'd54; b = 8'd254;  #10 
a = 8'd54; b = 8'd255;  #10 
a = 8'd55; b = 8'd0;  #10 
a = 8'd55; b = 8'd1;  #10 
a = 8'd55; b = 8'd2;  #10 
a = 8'd55; b = 8'd3;  #10 
a = 8'd55; b = 8'd4;  #10 
a = 8'd55; b = 8'd5;  #10 
a = 8'd55; b = 8'd6;  #10 
a = 8'd55; b = 8'd7;  #10 
a = 8'd55; b = 8'd8;  #10 
a = 8'd55; b = 8'd9;  #10 
a = 8'd55; b = 8'd10;  #10 
a = 8'd55; b = 8'd11;  #10 
a = 8'd55; b = 8'd12;  #10 
a = 8'd55; b = 8'd13;  #10 
a = 8'd55; b = 8'd14;  #10 
a = 8'd55; b = 8'd15;  #10 
a = 8'd55; b = 8'd16;  #10 
a = 8'd55; b = 8'd17;  #10 
a = 8'd55; b = 8'd18;  #10 
a = 8'd55; b = 8'd19;  #10 
a = 8'd55; b = 8'd20;  #10 
a = 8'd55; b = 8'd21;  #10 
a = 8'd55; b = 8'd22;  #10 
a = 8'd55; b = 8'd23;  #10 
a = 8'd55; b = 8'd24;  #10 
a = 8'd55; b = 8'd25;  #10 
a = 8'd55; b = 8'd26;  #10 
a = 8'd55; b = 8'd27;  #10 
a = 8'd55; b = 8'd28;  #10 
a = 8'd55; b = 8'd29;  #10 
a = 8'd55; b = 8'd30;  #10 
a = 8'd55; b = 8'd31;  #10 
a = 8'd55; b = 8'd32;  #10 
a = 8'd55; b = 8'd33;  #10 
a = 8'd55; b = 8'd34;  #10 
a = 8'd55; b = 8'd35;  #10 
a = 8'd55; b = 8'd36;  #10 
a = 8'd55; b = 8'd37;  #10 
a = 8'd55; b = 8'd38;  #10 
a = 8'd55; b = 8'd39;  #10 
a = 8'd55; b = 8'd40;  #10 
a = 8'd55; b = 8'd41;  #10 
a = 8'd55; b = 8'd42;  #10 
a = 8'd55; b = 8'd43;  #10 
a = 8'd55; b = 8'd44;  #10 
a = 8'd55; b = 8'd45;  #10 
a = 8'd55; b = 8'd46;  #10 
a = 8'd55; b = 8'd47;  #10 
a = 8'd55; b = 8'd48;  #10 
a = 8'd55; b = 8'd49;  #10 
a = 8'd55; b = 8'd50;  #10 
a = 8'd55; b = 8'd51;  #10 
a = 8'd55; b = 8'd52;  #10 
a = 8'd55; b = 8'd53;  #10 
a = 8'd55; b = 8'd54;  #10 
a = 8'd55; b = 8'd55;  #10 
a = 8'd55; b = 8'd56;  #10 
a = 8'd55; b = 8'd57;  #10 
a = 8'd55; b = 8'd58;  #10 
a = 8'd55; b = 8'd59;  #10 
a = 8'd55; b = 8'd60;  #10 
a = 8'd55; b = 8'd61;  #10 
a = 8'd55; b = 8'd62;  #10 
a = 8'd55; b = 8'd63;  #10 
a = 8'd55; b = 8'd64;  #10 
a = 8'd55; b = 8'd65;  #10 
a = 8'd55; b = 8'd66;  #10 
a = 8'd55; b = 8'd67;  #10 
a = 8'd55; b = 8'd68;  #10 
a = 8'd55; b = 8'd69;  #10 
a = 8'd55; b = 8'd70;  #10 
a = 8'd55; b = 8'd71;  #10 
a = 8'd55; b = 8'd72;  #10 
a = 8'd55; b = 8'd73;  #10 
a = 8'd55; b = 8'd74;  #10 
a = 8'd55; b = 8'd75;  #10 
a = 8'd55; b = 8'd76;  #10 
a = 8'd55; b = 8'd77;  #10 
a = 8'd55; b = 8'd78;  #10 
a = 8'd55; b = 8'd79;  #10 
a = 8'd55; b = 8'd80;  #10 
a = 8'd55; b = 8'd81;  #10 
a = 8'd55; b = 8'd82;  #10 
a = 8'd55; b = 8'd83;  #10 
a = 8'd55; b = 8'd84;  #10 
a = 8'd55; b = 8'd85;  #10 
a = 8'd55; b = 8'd86;  #10 
a = 8'd55; b = 8'd87;  #10 
a = 8'd55; b = 8'd88;  #10 
a = 8'd55; b = 8'd89;  #10 
a = 8'd55; b = 8'd90;  #10 
a = 8'd55; b = 8'd91;  #10 
a = 8'd55; b = 8'd92;  #10 
a = 8'd55; b = 8'd93;  #10 
a = 8'd55; b = 8'd94;  #10 
a = 8'd55; b = 8'd95;  #10 
a = 8'd55; b = 8'd96;  #10 
a = 8'd55; b = 8'd97;  #10 
a = 8'd55; b = 8'd98;  #10 
a = 8'd55; b = 8'd99;  #10 
a = 8'd55; b = 8'd100;  #10 
a = 8'd55; b = 8'd101;  #10 
a = 8'd55; b = 8'd102;  #10 
a = 8'd55; b = 8'd103;  #10 
a = 8'd55; b = 8'd104;  #10 
a = 8'd55; b = 8'd105;  #10 
a = 8'd55; b = 8'd106;  #10 
a = 8'd55; b = 8'd107;  #10 
a = 8'd55; b = 8'd108;  #10 
a = 8'd55; b = 8'd109;  #10 
a = 8'd55; b = 8'd110;  #10 
a = 8'd55; b = 8'd111;  #10 
a = 8'd55; b = 8'd112;  #10 
a = 8'd55; b = 8'd113;  #10 
a = 8'd55; b = 8'd114;  #10 
a = 8'd55; b = 8'd115;  #10 
a = 8'd55; b = 8'd116;  #10 
a = 8'd55; b = 8'd117;  #10 
a = 8'd55; b = 8'd118;  #10 
a = 8'd55; b = 8'd119;  #10 
a = 8'd55; b = 8'd120;  #10 
a = 8'd55; b = 8'd121;  #10 
a = 8'd55; b = 8'd122;  #10 
a = 8'd55; b = 8'd123;  #10 
a = 8'd55; b = 8'd124;  #10 
a = 8'd55; b = 8'd125;  #10 
a = 8'd55; b = 8'd126;  #10 
a = 8'd55; b = 8'd127;  #10 
a = 8'd55; b = 8'd128;  #10 
a = 8'd55; b = 8'd129;  #10 
a = 8'd55; b = 8'd130;  #10 
a = 8'd55; b = 8'd131;  #10 
a = 8'd55; b = 8'd132;  #10 
a = 8'd55; b = 8'd133;  #10 
a = 8'd55; b = 8'd134;  #10 
a = 8'd55; b = 8'd135;  #10 
a = 8'd55; b = 8'd136;  #10 
a = 8'd55; b = 8'd137;  #10 
a = 8'd55; b = 8'd138;  #10 
a = 8'd55; b = 8'd139;  #10 
a = 8'd55; b = 8'd140;  #10 
a = 8'd55; b = 8'd141;  #10 
a = 8'd55; b = 8'd142;  #10 
a = 8'd55; b = 8'd143;  #10 
a = 8'd55; b = 8'd144;  #10 
a = 8'd55; b = 8'd145;  #10 
a = 8'd55; b = 8'd146;  #10 
a = 8'd55; b = 8'd147;  #10 
a = 8'd55; b = 8'd148;  #10 
a = 8'd55; b = 8'd149;  #10 
a = 8'd55; b = 8'd150;  #10 
a = 8'd55; b = 8'd151;  #10 
a = 8'd55; b = 8'd152;  #10 
a = 8'd55; b = 8'd153;  #10 
a = 8'd55; b = 8'd154;  #10 
a = 8'd55; b = 8'd155;  #10 
a = 8'd55; b = 8'd156;  #10 
a = 8'd55; b = 8'd157;  #10 
a = 8'd55; b = 8'd158;  #10 
a = 8'd55; b = 8'd159;  #10 
a = 8'd55; b = 8'd160;  #10 
a = 8'd55; b = 8'd161;  #10 
a = 8'd55; b = 8'd162;  #10 
a = 8'd55; b = 8'd163;  #10 
a = 8'd55; b = 8'd164;  #10 
a = 8'd55; b = 8'd165;  #10 
a = 8'd55; b = 8'd166;  #10 
a = 8'd55; b = 8'd167;  #10 
a = 8'd55; b = 8'd168;  #10 
a = 8'd55; b = 8'd169;  #10 
a = 8'd55; b = 8'd170;  #10 
a = 8'd55; b = 8'd171;  #10 
a = 8'd55; b = 8'd172;  #10 
a = 8'd55; b = 8'd173;  #10 
a = 8'd55; b = 8'd174;  #10 
a = 8'd55; b = 8'd175;  #10 
a = 8'd55; b = 8'd176;  #10 
a = 8'd55; b = 8'd177;  #10 
a = 8'd55; b = 8'd178;  #10 
a = 8'd55; b = 8'd179;  #10 
a = 8'd55; b = 8'd180;  #10 
a = 8'd55; b = 8'd181;  #10 
a = 8'd55; b = 8'd182;  #10 
a = 8'd55; b = 8'd183;  #10 
a = 8'd55; b = 8'd184;  #10 
a = 8'd55; b = 8'd185;  #10 
a = 8'd55; b = 8'd186;  #10 
a = 8'd55; b = 8'd187;  #10 
a = 8'd55; b = 8'd188;  #10 
a = 8'd55; b = 8'd189;  #10 
a = 8'd55; b = 8'd190;  #10 
a = 8'd55; b = 8'd191;  #10 
a = 8'd55; b = 8'd192;  #10 
a = 8'd55; b = 8'd193;  #10 
a = 8'd55; b = 8'd194;  #10 
a = 8'd55; b = 8'd195;  #10 
a = 8'd55; b = 8'd196;  #10 
a = 8'd55; b = 8'd197;  #10 
a = 8'd55; b = 8'd198;  #10 
a = 8'd55; b = 8'd199;  #10 
a = 8'd55; b = 8'd200;  #10 
a = 8'd55; b = 8'd201;  #10 
a = 8'd55; b = 8'd202;  #10 
a = 8'd55; b = 8'd203;  #10 
a = 8'd55; b = 8'd204;  #10 
a = 8'd55; b = 8'd205;  #10 
a = 8'd55; b = 8'd206;  #10 
a = 8'd55; b = 8'd207;  #10 
a = 8'd55; b = 8'd208;  #10 
a = 8'd55; b = 8'd209;  #10 
a = 8'd55; b = 8'd210;  #10 
a = 8'd55; b = 8'd211;  #10 
a = 8'd55; b = 8'd212;  #10 
a = 8'd55; b = 8'd213;  #10 
a = 8'd55; b = 8'd214;  #10 
a = 8'd55; b = 8'd215;  #10 
a = 8'd55; b = 8'd216;  #10 
a = 8'd55; b = 8'd217;  #10 
a = 8'd55; b = 8'd218;  #10 
a = 8'd55; b = 8'd219;  #10 
a = 8'd55; b = 8'd220;  #10 
a = 8'd55; b = 8'd221;  #10 
a = 8'd55; b = 8'd222;  #10 
a = 8'd55; b = 8'd223;  #10 
a = 8'd55; b = 8'd224;  #10 
a = 8'd55; b = 8'd225;  #10 
a = 8'd55; b = 8'd226;  #10 
a = 8'd55; b = 8'd227;  #10 
a = 8'd55; b = 8'd228;  #10 
a = 8'd55; b = 8'd229;  #10 
a = 8'd55; b = 8'd230;  #10 
a = 8'd55; b = 8'd231;  #10 
a = 8'd55; b = 8'd232;  #10 
a = 8'd55; b = 8'd233;  #10 
a = 8'd55; b = 8'd234;  #10 
a = 8'd55; b = 8'd235;  #10 
a = 8'd55; b = 8'd236;  #10 
a = 8'd55; b = 8'd237;  #10 
a = 8'd55; b = 8'd238;  #10 
a = 8'd55; b = 8'd239;  #10 
a = 8'd55; b = 8'd240;  #10 
a = 8'd55; b = 8'd241;  #10 
a = 8'd55; b = 8'd242;  #10 
a = 8'd55; b = 8'd243;  #10 
a = 8'd55; b = 8'd244;  #10 
a = 8'd55; b = 8'd245;  #10 
a = 8'd55; b = 8'd246;  #10 
a = 8'd55; b = 8'd247;  #10 
a = 8'd55; b = 8'd248;  #10 
a = 8'd55; b = 8'd249;  #10 
a = 8'd55; b = 8'd250;  #10 
a = 8'd55; b = 8'd251;  #10 
a = 8'd55; b = 8'd252;  #10 
a = 8'd55; b = 8'd253;  #10 
a = 8'd55; b = 8'd254;  #10 
a = 8'd55; b = 8'd255;  #10 
a = 8'd56; b = 8'd0;  #10 
a = 8'd56; b = 8'd1;  #10 
a = 8'd56; b = 8'd2;  #10 
a = 8'd56; b = 8'd3;  #10 
a = 8'd56; b = 8'd4;  #10 
a = 8'd56; b = 8'd5;  #10 
a = 8'd56; b = 8'd6;  #10 
a = 8'd56; b = 8'd7;  #10 
a = 8'd56; b = 8'd8;  #10 
a = 8'd56; b = 8'd9;  #10 
a = 8'd56; b = 8'd10;  #10 
a = 8'd56; b = 8'd11;  #10 
a = 8'd56; b = 8'd12;  #10 
a = 8'd56; b = 8'd13;  #10 
a = 8'd56; b = 8'd14;  #10 
a = 8'd56; b = 8'd15;  #10 
a = 8'd56; b = 8'd16;  #10 
a = 8'd56; b = 8'd17;  #10 
a = 8'd56; b = 8'd18;  #10 
a = 8'd56; b = 8'd19;  #10 
a = 8'd56; b = 8'd20;  #10 
a = 8'd56; b = 8'd21;  #10 
a = 8'd56; b = 8'd22;  #10 
a = 8'd56; b = 8'd23;  #10 
a = 8'd56; b = 8'd24;  #10 
a = 8'd56; b = 8'd25;  #10 
a = 8'd56; b = 8'd26;  #10 
a = 8'd56; b = 8'd27;  #10 
a = 8'd56; b = 8'd28;  #10 
a = 8'd56; b = 8'd29;  #10 
a = 8'd56; b = 8'd30;  #10 
a = 8'd56; b = 8'd31;  #10 
a = 8'd56; b = 8'd32;  #10 
a = 8'd56; b = 8'd33;  #10 
a = 8'd56; b = 8'd34;  #10 
a = 8'd56; b = 8'd35;  #10 
a = 8'd56; b = 8'd36;  #10 
a = 8'd56; b = 8'd37;  #10 
a = 8'd56; b = 8'd38;  #10 
a = 8'd56; b = 8'd39;  #10 
a = 8'd56; b = 8'd40;  #10 
a = 8'd56; b = 8'd41;  #10 
a = 8'd56; b = 8'd42;  #10 
a = 8'd56; b = 8'd43;  #10 
a = 8'd56; b = 8'd44;  #10 
a = 8'd56; b = 8'd45;  #10 
a = 8'd56; b = 8'd46;  #10 
a = 8'd56; b = 8'd47;  #10 
a = 8'd56; b = 8'd48;  #10 
a = 8'd56; b = 8'd49;  #10 
a = 8'd56; b = 8'd50;  #10 
a = 8'd56; b = 8'd51;  #10 
a = 8'd56; b = 8'd52;  #10 
a = 8'd56; b = 8'd53;  #10 
a = 8'd56; b = 8'd54;  #10 
a = 8'd56; b = 8'd55;  #10 
a = 8'd56; b = 8'd56;  #10 
a = 8'd56; b = 8'd57;  #10 
a = 8'd56; b = 8'd58;  #10 
a = 8'd56; b = 8'd59;  #10 
a = 8'd56; b = 8'd60;  #10 
a = 8'd56; b = 8'd61;  #10 
a = 8'd56; b = 8'd62;  #10 
a = 8'd56; b = 8'd63;  #10 
a = 8'd56; b = 8'd64;  #10 
a = 8'd56; b = 8'd65;  #10 
a = 8'd56; b = 8'd66;  #10 
a = 8'd56; b = 8'd67;  #10 
a = 8'd56; b = 8'd68;  #10 
a = 8'd56; b = 8'd69;  #10 
a = 8'd56; b = 8'd70;  #10 
a = 8'd56; b = 8'd71;  #10 
a = 8'd56; b = 8'd72;  #10 
a = 8'd56; b = 8'd73;  #10 
a = 8'd56; b = 8'd74;  #10 
a = 8'd56; b = 8'd75;  #10 
a = 8'd56; b = 8'd76;  #10 
a = 8'd56; b = 8'd77;  #10 
a = 8'd56; b = 8'd78;  #10 
a = 8'd56; b = 8'd79;  #10 
a = 8'd56; b = 8'd80;  #10 
a = 8'd56; b = 8'd81;  #10 
a = 8'd56; b = 8'd82;  #10 
a = 8'd56; b = 8'd83;  #10 
a = 8'd56; b = 8'd84;  #10 
a = 8'd56; b = 8'd85;  #10 
a = 8'd56; b = 8'd86;  #10 
a = 8'd56; b = 8'd87;  #10 
a = 8'd56; b = 8'd88;  #10 
a = 8'd56; b = 8'd89;  #10 
a = 8'd56; b = 8'd90;  #10 
a = 8'd56; b = 8'd91;  #10 
a = 8'd56; b = 8'd92;  #10 
a = 8'd56; b = 8'd93;  #10 
a = 8'd56; b = 8'd94;  #10 
a = 8'd56; b = 8'd95;  #10 
a = 8'd56; b = 8'd96;  #10 
a = 8'd56; b = 8'd97;  #10 
a = 8'd56; b = 8'd98;  #10 
a = 8'd56; b = 8'd99;  #10 
a = 8'd56; b = 8'd100;  #10 
a = 8'd56; b = 8'd101;  #10 
a = 8'd56; b = 8'd102;  #10 
a = 8'd56; b = 8'd103;  #10 
a = 8'd56; b = 8'd104;  #10 
a = 8'd56; b = 8'd105;  #10 
a = 8'd56; b = 8'd106;  #10 
a = 8'd56; b = 8'd107;  #10 
a = 8'd56; b = 8'd108;  #10 
a = 8'd56; b = 8'd109;  #10 
a = 8'd56; b = 8'd110;  #10 
a = 8'd56; b = 8'd111;  #10 
a = 8'd56; b = 8'd112;  #10 
a = 8'd56; b = 8'd113;  #10 
a = 8'd56; b = 8'd114;  #10 
a = 8'd56; b = 8'd115;  #10 
a = 8'd56; b = 8'd116;  #10 
a = 8'd56; b = 8'd117;  #10 
a = 8'd56; b = 8'd118;  #10 
a = 8'd56; b = 8'd119;  #10 
a = 8'd56; b = 8'd120;  #10 
a = 8'd56; b = 8'd121;  #10 
a = 8'd56; b = 8'd122;  #10 
a = 8'd56; b = 8'd123;  #10 
a = 8'd56; b = 8'd124;  #10 
a = 8'd56; b = 8'd125;  #10 
a = 8'd56; b = 8'd126;  #10 
a = 8'd56; b = 8'd127;  #10 
a = 8'd56; b = 8'd128;  #10 
a = 8'd56; b = 8'd129;  #10 
a = 8'd56; b = 8'd130;  #10 
a = 8'd56; b = 8'd131;  #10 
a = 8'd56; b = 8'd132;  #10 
a = 8'd56; b = 8'd133;  #10 
a = 8'd56; b = 8'd134;  #10 
a = 8'd56; b = 8'd135;  #10 
a = 8'd56; b = 8'd136;  #10 
a = 8'd56; b = 8'd137;  #10 
a = 8'd56; b = 8'd138;  #10 
a = 8'd56; b = 8'd139;  #10 
a = 8'd56; b = 8'd140;  #10 
a = 8'd56; b = 8'd141;  #10 
a = 8'd56; b = 8'd142;  #10 
a = 8'd56; b = 8'd143;  #10 
a = 8'd56; b = 8'd144;  #10 
a = 8'd56; b = 8'd145;  #10 
a = 8'd56; b = 8'd146;  #10 
a = 8'd56; b = 8'd147;  #10 
a = 8'd56; b = 8'd148;  #10 
a = 8'd56; b = 8'd149;  #10 
a = 8'd56; b = 8'd150;  #10 
a = 8'd56; b = 8'd151;  #10 
a = 8'd56; b = 8'd152;  #10 
a = 8'd56; b = 8'd153;  #10 
a = 8'd56; b = 8'd154;  #10 
a = 8'd56; b = 8'd155;  #10 
a = 8'd56; b = 8'd156;  #10 
a = 8'd56; b = 8'd157;  #10 
a = 8'd56; b = 8'd158;  #10 
a = 8'd56; b = 8'd159;  #10 
a = 8'd56; b = 8'd160;  #10 
a = 8'd56; b = 8'd161;  #10 
a = 8'd56; b = 8'd162;  #10 
a = 8'd56; b = 8'd163;  #10 
a = 8'd56; b = 8'd164;  #10 
a = 8'd56; b = 8'd165;  #10 
a = 8'd56; b = 8'd166;  #10 
a = 8'd56; b = 8'd167;  #10 
a = 8'd56; b = 8'd168;  #10 
a = 8'd56; b = 8'd169;  #10 
a = 8'd56; b = 8'd170;  #10 
a = 8'd56; b = 8'd171;  #10 
a = 8'd56; b = 8'd172;  #10 
a = 8'd56; b = 8'd173;  #10 
a = 8'd56; b = 8'd174;  #10 
a = 8'd56; b = 8'd175;  #10 
a = 8'd56; b = 8'd176;  #10 
a = 8'd56; b = 8'd177;  #10 
a = 8'd56; b = 8'd178;  #10 
a = 8'd56; b = 8'd179;  #10 
a = 8'd56; b = 8'd180;  #10 
a = 8'd56; b = 8'd181;  #10 
a = 8'd56; b = 8'd182;  #10 
a = 8'd56; b = 8'd183;  #10 
a = 8'd56; b = 8'd184;  #10 
a = 8'd56; b = 8'd185;  #10 
a = 8'd56; b = 8'd186;  #10 
a = 8'd56; b = 8'd187;  #10 
a = 8'd56; b = 8'd188;  #10 
a = 8'd56; b = 8'd189;  #10 
a = 8'd56; b = 8'd190;  #10 
a = 8'd56; b = 8'd191;  #10 
a = 8'd56; b = 8'd192;  #10 
a = 8'd56; b = 8'd193;  #10 
a = 8'd56; b = 8'd194;  #10 
a = 8'd56; b = 8'd195;  #10 
a = 8'd56; b = 8'd196;  #10 
a = 8'd56; b = 8'd197;  #10 
a = 8'd56; b = 8'd198;  #10 
a = 8'd56; b = 8'd199;  #10 
a = 8'd56; b = 8'd200;  #10 
a = 8'd56; b = 8'd201;  #10 
a = 8'd56; b = 8'd202;  #10 
a = 8'd56; b = 8'd203;  #10 
a = 8'd56; b = 8'd204;  #10 
a = 8'd56; b = 8'd205;  #10 
a = 8'd56; b = 8'd206;  #10 
a = 8'd56; b = 8'd207;  #10 
a = 8'd56; b = 8'd208;  #10 
a = 8'd56; b = 8'd209;  #10 
a = 8'd56; b = 8'd210;  #10 
a = 8'd56; b = 8'd211;  #10 
a = 8'd56; b = 8'd212;  #10 
a = 8'd56; b = 8'd213;  #10 
a = 8'd56; b = 8'd214;  #10 
a = 8'd56; b = 8'd215;  #10 
a = 8'd56; b = 8'd216;  #10 
a = 8'd56; b = 8'd217;  #10 
a = 8'd56; b = 8'd218;  #10 
a = 8'd56; b = 8'd219;  #10 
a = 8'd56; b = 8'd220;  #10 
a = 8'd56; b = 8'd221;  #10 
a = 8'd56; b = 8'd222;  #10 
a = 8'd56; b = 8'd223;  #10 
a = 8'd56; b = 8'd224;  #10 
a = 8'd56; b = 8'd225;  #10 
a = 8'd56; b = 8'd226;  #10 
a = 8'd56; b = 8'd227;  #10 
a = 8'd56; b = 8'd228;  #10 
a = 8'd56; b = 8'd229;  #10 
a = 8'd56; b = 8'd230;  #10 
a = 8'd56; b = 8'd231;  #10 
a = 8'd56; b = 8'd232;  #10 
a = 8'd56; b = 8'd233;  #10 
a = 8'd56; b = 8'd234;  #10 
a = 8'd56; b = 8'd235;  #10 
a = 8'd56; b = 8'd236;  #10 
a = 8'd56; b = 8'd237;  #10 
a = 8'd56; b = 8'd238;  #10 
a = 8'd56; b = 8'd239;  #10 
a = 8'd56; b = 8'd240;  #10 
a = 8'd56; b = 8'd241;  #10 
a = 8'd56; b = 8'd242;  #10 
a = 8'd56; b = 8'd243;  #10 
a = 8'd56; b = 8'd244;  #10 
a = 8'd56; b = 8'd245;  #10 
a = 8'd56; b = 8'd246;  #10 
a = 8'd56; b = 8'd247;  #10 
a = 8'd56; b = 8'd248;  #10 
a = 8'd56; b = 8'd249;  #10 
a = 8'd56; b = 8'd250;  #10 
a = 8'd56; b = 8'd251;  #10 
a = 8'd56; b = 8'd252;  #10 
a = 8'd56; b = 8'd253;  #10 
a = 8'd56; b = 8'd254;  #10 
a = 8'd56; b = 8'd255;  #10 
a = 8'd57; b = 8'd0;  #10 
a = 8'd57; b = 8'd1;  #10 
a = 8'd57; b = 8'd2;  #10 
a = 8'd57; b = 8'd3;  #10 
a = 8'd57; b = 8'd4;  #10 
a = 8'd57; b = 8'd5;  #10 
a = 8'd57; b = 8'd6;  #10 
a = 8'd57; b = 8'd7;  #10 
a = 8'd57; b = 8'd8;  #10 
a = 8'd57; b = 8'd9;  #10 
a = 8'd57; b = 8'd10;  #10 
a = 8'd57; b = 8'd11;  #10 
a = 8'd57; b = 8'd12;  #10 
a = 8'd57; b = 8'd13;  #10 
a = 8'd57; b = 8'd14;  #10 
a = 8'd57; b = 8'd15;  #10 
a = 8'd57; b = 8'd16;  #10 
a = 8'd57; b = 8'd17;  #10 
a = 8'd57; b = 8'd18;  #10 
a = 8'd57; b = 8'd19;  #10 
a = 8'd57; b = 8'd20;  #10 
a = 8'd57; b = 8'd21;  #10 
a = 8'd57; b = 8'd22;  #10 
a = 8'd57; b = 8'd23;  #10 
a = 8'd57; b = 8'd24;  #10 
a = 8'd57; b = 8'd25;  #10 
a = 8'd57; b = 8'd26;  #10 
a = 8'd57; b = 8'd27;  #10 
a = 8'd57; b = 8'd28;  #10 
a = 8'd57; b = 8'd29;  #10 
a = 8'd57; b = 8'd30;  #10 
a = 8'd57; b = 8'd31;  #10 
a = 8'd57; b = 8'd32;  #10 
a = 8'd57; b = 8'd33;  #10 
a = 8'd57; b = 8'd34;  #10 
a = 8'd57; b = 8'd35;  #10 
a = 8'd57; b = 8'd36;  #10 
a = 8'd57; b = 8'd37;  #10 
a = 8'd57; b = 8'd38;  #10 
a = 8'd57; b = 8'd39;  #10 
a = 8'd57; b = 8'd40;  #10 
a = 8'd57; b = 8'd41;  #10 
a = 8'd57; b = 8'd42;  #10 
a = 8'd57; b = 8'd43;  #10 
a = 8'd57; b = 8'd44;  #10 
a = 8'd57; b = 8'd45;  #10 
a = 8'd57; b = 8'd46;  #10 
a = 8'd57; b = 8'd47;  #10 
a = 8'd57; b = 8'd48;  #10 
a = 8'd57; b = 8'd49;  #10 
a = 8'd57; b = 8'd50;  #10 
a = 8'd57; b = 8'd51;  #10 
a = 8'd57; b = 8'd52;  #10 
a = 8'd57; b = 8'd53;  #10 
a = 8'd57; b = 8'd54;  #10 
a = 8'd57; b = 8'd55;  #10 
a = 8'd57; b = 8'd56;  #10 
a = 8'd57; b = 8'd57;  #10 
a = 8'd57; b = 8'd58;  #10 
a = 8'd57; b = 8'd59;  #10 
a = 8'd57; b = 8'd60;  #10 
a = 8'd57; b = 8'd61;  #10 
a = 8'd57; b = 8'd62;  #10 
a = 8'd57; b = 8'd63;  #10 
a = 8'd57; b = 8'd64;  #10 
a = 8'd57; b = 8'd65;  #10 
a = 8'd57; b = 8'd66;  #10 
a = 8'd57; b = 8'd67;  #10 
a = 8'd57; b = 8'd68;  #10 
a = 8'd57; b = 8'd69;  #10 
a = 8'd57; b = 8'd70;  #10 
a = 8'd57; b = 8'd71;  #10 
a = 8'd57; b = 8'd72;  #10 
a = 8'd57; b = 8'd73;  #10 
a = 8'd57; b = 8'd74;  #10 
a = 8'd57; b = 8'd75;  #10 
a = 8'd57; b = 8'd76;  #10 
a = 8'd57; b = 8'd77;  #10 
a = 8'd57; b = 8'd78;  #10 
a = 8'd57; b = 8'd79;  #10 
a = 8'd57; b = 8'd80;  #10 
a = 8'd57; b = 8'd81;  #10 
a = 8'd57; b = 8'd82;  #10 
a = 8'd57; b = 8'd83;  #10 
a = 8'd57; b = 8'd84;  #10 
a = 8'd57; b = 8'd85;  #10 
a = 8'd57; b = 8'd86;  #10 
a = 8'd57; b = 8'd87;  #10 
a = 8'd57; b = 8'd88;  #10 
a = 8'd57; b = 8'd89;  #10 
a = 8'd57; b = 8'd90;  #10 
a = 8'd57; b = 8'd91;  #10 
a = 8'd57; b = 8'd92;  #10 
a = 8'd57; b = 8'd93;  #10 
a = 8'd57; b = 8'd94;  #10 
a = 8'd57; b = 8'd95;  #10 
a = 8'd57; b = 8'd96;  #10 
a = 8'd57; b = 8'd97;  #10 
a = 8'd57; b = 8'd98;  #10 
a = 8'd57; b = 8'd99;  #10 
a = 8'd57; b = 8'd100;  #10 
a = 8'd57; b = 8'd101;  #10 
a = 8'd57; b = 8'd102;  #10 
a = 8'd57; b = 8'd103;  #10 
a = 8'd57; b = 8'd104;  #10 
a = 8'd57; b = 8'd105;  #10 
a = 8'd57; b = 8'd106;  #10 
a = 8'd57; b = 8'd107;  #10 
a = 8'd57; b = 8'd108;  #10 
a = 8'd57; b = 8'd109;  #10 
a = 8'd57; b = 8'd110;  #10 
a = 8'd57; b = 8'd111;  #10 
a = 8'd57; b = 8'd112;  #10 
a = 8'd57; b = 8'd113;  #10 
a = 8'd57; b = 8'd114;  #10 
a = 8'd57; b = 8'd115;  #10 
a = 8'd57; b = 8'd116;  #10 
a = 8'd57; b = 8'd117;  #10 
a = 8'd57; b = 8'd118;  #10 
a = 8'd57; b = 8'd119;  #10 
a = 8'd57; b = 8'd120;  #10 
a = 8'd57; b = 8'd121;  #10 
a = 8'd57; b = 8'd122;  #10 
a = 8'd57; b = 8'd123;  #10 
a = 8'd57; b = 8'd124;  #10 
a = 8'd57; b = 8'd125;  #10 
a = 8'd57; b = 8'd126;  #10 
a = 8'd57; b = 8'd127;  #10 
a = 8'd57; b = 8'd128;  #10 
a = 8'd57; b = 8'd129;  #10 
a = 8'd57; b = 8'd130;  #10 
a = 8'd57; b = 8'd131;  #10 
a = 8'd57; b = 8'd132;  #10 
a = 8'd57; b = 8'd133;  #10 
a = 8'd57; b = 8'd134;  #10 
a = 8'd57; b = 8'd135;  #10 
a = 8'd57; b = 8'd136;  #10 
a = 8'd57; b = 8'd137;  #10 
a = 8'd57; b = 8'd138;  #10 
a = 8'd57; b = 8'd139;  #10 
a = 8'd57; b = 8'd140;  #10 
a = 8'd57; b = 8'd141;  #10 
a = 8'd57; b = 8'd142;  #10 
a = 8'd57; b = 8'd143;  #10 
a = 8'd57; b = 8'd144;  #10 
a = 8'd57; b = 8'd145;  #10 
a = 8'd57; b = 8'd146;  #10 
a = 8'd57; b = 8'd147;  #10 
a = 8'd57; b = 8'd148;  #10 
a = 8'd57; b = 8'd149;  #10 
a = 8'd57; b = 8'd150;  #10 
a = 8'd57; b = 8'd151;  #10 
a = 8'd57; b = 8'd152;  #10 
a = 8'd57; b = 8'd153;  #10 
a = 8'd57; b = 8'd154;  #10 
a = 8'd57; b = 8'd155;  #10 
a = 8'd57; b = 8'd156;  #10 
a = 8'd57; b = 8'd157;  #10 
a = 8'd57; b = 8'd158;  #10 
a = 8'd57; b = 8'd159;  #10 
a = 8'd57; b = 8'd160;  #10 
a = 8'd57; b = 8'd161;  #10 
a = 8'd57; b = 8'd162;  #10 
a = 8'd57; b = 8'd163;  #10 
a = 8'd57; b = 8'd164;  #10 
a = 8'd57; b = 8'd165;  #10 
a = 8'd57; b = 8'd166;  #10 
a = 8'd57; b = 8'd167;  #10 
a = 8'd57; b = 8'd168;  #10 
a = 8'd57; b = 8'd169;  #10 
a = 8'd57; b = 8'd170;  #10 
a = 8'd57; b = 8'd171;  #10 
a = 8'd57; b = 8'd172;  #10 
a = 8'd57; b = 8'd173;  #10 
a = 8'd57; b = 8'd174;  #10 
a = 8'd57; b = 8'd175;  #10 
a = 8'd57; b = 8'd176;  #10 
a = 8'd57; b = 8'd177;  #10 
a = 8'd57; b = 8'd178;  #10 
a = 8'd57; b = 8'd179;  #10 
a = 8'd57; b = 8'd180;  #10 
a = 8'd57; b = 8'd181;  #10 
a = 8'd57; b = 8'd182;  #10 
a = 8'd57; b = 8'd183;  #10 
a = 8'd57; b = 8'd184;  #10 
a = 8'd57; b = 8'd185;  #10 
a = 8'd57; b = 8'd186;  #10 
a = 8'd57; b = 8'd187;  #10 
a = 8'd57; b = 8'd188;  #10 
a = 8'd57; b = 8'd189;  #10 
a = 8'd57; b = 8'd190;  #10 
a = 8'd57; b = 8'd191;  #10 
a = 8'd57; b = 8'd192;  #10 
a = 8'd57; b = 8'd193;  #10 
a = 8'd57; b = 8'd194;  #10 
a = 8'd57; b = 8'd195;  #10 
a = 8'd57; b = 8'd196;  #10 
a = 8'd57; b = 8'd197;  #10 
a = 8'd57; b = 8'd198;  #10 
a = 8'd57; b = 8'd199;  #10 
a = 8'd57; b = 8'd200;  #10 
a = 8'd57; b = 8'd201;  #10 
a = 8'd57; b = 8'd202;  #10 
a = 8'd57; b = 8'd203;  #10 
a = 8'd57; b = 8'd204;  #10 
a = 8'd57; b = 8'd205;  #10 
a = 8'd57; b = 8'd206;  #10 
a = 8'd57; b = 8'd207;  #10 
a = 8'd57; b = 8'd208;  #10 
a = 8'd57; b = 8'd209;  #10 
a = 8'd57; b = 8'd210;  #10 
a = 8'd57; b = 8'd211;  #10 
a = 8'd57; b = 8'd212;  #10 
a = 8'd57; b = 8'd213;  #10 
a = 8'd57; b = 8'd214;  #10 
a = 8'd57; b = 8'd215;  #10 
a = 8'd57; b = 8'd216;  #10 
a = 8'd57; b = 8'd217;  #10 
a = 8'd57; b = 8'd218;  #10 
a = 8'd57; b = 8'd219;  #10 
a = 8'd57; b = 8'd220;  #10 
a = 8'd57; b = 8'd221;  #10 
a = 8'd57; b = 8'd222;  #10 
a = 8'd57; b = 8'd223;  #10 
a = 8'd57; b = 8'd224;  #10 
a = 8'd57; b = 8'd225;  #10 
a = 8'd57; b = 8'd226;  #10 
a = 8'd57; b = 8'd227;  #10 
a = 8'd57; b = 8'd228;  #10 
a = 8'd57; b = 8'd229;  #10 
a = 8'd57; b = 8'd230;  #10 
a = 8'd57; b = 8'd231;  #10 
a = 8'd57; b = 8'd232;  #10 
a = 8'd57; b = 8'd233;  #10 
a = 8'd57; b = 8'd234;  #10 
a = 8'd57; b = 8'd235;  #10 
a = 8'd57; b = 8'd236;  #10 
a = 8'd57; b = 8'd237;  #10 
a = 8'd57; b = 8'd238;  #10 
a = 8'd57; b = 8'd239;  #10 
a = 8'd57; b = 8'd240;  #10 
a = 8'd57; b = 8'd241;  #10 
a = 8'd57; b = 8'd242;  #10 
a = 8'd57; b = 8'd243;  #10 
a = 8'd57; b = 8'd244;  #10 
a = 8'd57; b = 8'd245;  #10 
a = 8'd57; b = 8'd246;  #10 
a = 8'd57; b = 8'd247;  #10 
a = 8'd57; b = 8'd248;  #10 
a = 8'd57; b = 8'd249;  #10 
a = 8'd57; b = 8'd250;  #10 
a = 8'd57; b = 8'd251;  #10 
a = 8'd57; b = 8'd252;  #10 
a = 8'd57; b = 8'd253;  #10 
a = 8'd57; b = 8'd254;  #10 
a = 8'd57; b = 8'd255;  #10 
a = 8'd58; b = 8'd0;  #10 
a = 8'd58; b = 8'd1;  #10 
a = 8'd58; b = 8'd2;  #10 
a = 8'd58; b = 8'd3;  #10 
a = 8'd58; b = 8'd4;  #10 
a = 8'd58; b = 8'd5;  #10 
a = 8'd58; b = 8'd6;  #10 
a = 8'd58; b = 8'd7;  #10 
a = 8'd58; b = 8'd8;  #10 
a = 8'd58; b = 8'd9;  #10 
a = 8'd58; b = 8'd10;  #10 
a = 8'd58; b = 8'd11;  #10 
a = 8'd58; b = 8'd12;  #10 
a = 8'd58; b = 8'd13;  #10 
a = 8'd58; b = 8'd14;  #10 
a = 8'd58; b = 8'd15;  #10 
a = 8'd58; b = 8'd16;  #10 
a = 8'd58; b = 8'd17;  #10 
a = 8'd58; b = 8'd18;  #10 
a = 8'd58; b = 8'd19;  #10 
a = 8'd58; b = 8'd20;  #10 
a = 8'd58; b = 8'd21;  #10 
a = 8'd58; b = 8'd22;  #10 
a = 8'd58; b = 8'd23;  #10 
a = 8'd58; b = 8'd24;  #10 
a = 8'd58; b = 8'd25;  #10 
a = 8'd58; b = 8'd26;  #10 
a = 8'd58; b = 8'd27;  #10 
a = 8'd58; b = 8'd28;  #10 
a = 8'd58; b = 8'd29;  #10 
a = 8'd58; b = 8'd30;  #10 
a = 8'd58; b = 8'd31;  #10 
a = 8'd58; b = 8'd32;  #10 
a = 8'd58; b = 8'd33;  #10 
a = 8'd58; b = 8'd34;  #10 
a = 8'd58; b = 8'd35;  #10 
a = 8'd58; b = 8'd36;  #10 
a = 8'd58; b = 8'd37;  #10 
a = 8'd58; b = 8'd38;  #10 
a = 8'd58; b = 8'd39;  #10 
a = 8'd58; b = 8'd40;  #10 
a = 8'd58; b = 8'd41;  #10 
a = 8'd58; b = 8'd42;  #10 
a = 8'd58; b = 8'd43;  #10 
a = 8'd58; b = 8'd44;  #10 
a = 8'd58; b = 8'd45;  #10 
a = 8'd58; b = 8'd46;  #10 
a = 8'd58; b = 8'd47;  #10 
a = 8'd58; b = 8'd48;  #10 
a = 8'd58; b = 8'd49;  #10 
a = 8'd58; b = 8'd50;  #10 
a = 8'd58; b = 8'd51;  #10 
a = 8'd58; b = 8'd52;  #10 
a = 8'd58; b = 8'd53;  #10 
a = 8'd58; b = 8'd54;  #10 
a = 8'd58; b = 8'd55;  #10 
a = 8'd58; b = 8'd56;  #10 
a = 8'd58; b = 8'd57;  #10 
a = 8'd58; b = 8'd58;  #10 
a = 8'd58; b = 8'd59;  #10 
a = 8'd58; b = 8'd60;  #10 
a = 8'd58; b = 8'd61;  #10 
a = 8'd58; b = 8'd62;  #10 
a = 8'd58; b = 8'd63;  #10 
a = 8'd58; b = 8'd64;  #10 
a = 8'd58; b = 8'd65;  #10 
a = 8'd58; b = 8'd66;  #10 
a = 8'd58; b = 8'd67;  #10 
a = 8'd58; b = 8'd68;  #10 
a = 8'd58; b = 8'd69;  #10 
a = 8'd58; b = 8'd70;  #10 
a = 8'd58; b = 8'd71;  #10 
a = 8'd58; b = 8'd72;  #10 
a = 8'd58; b = 8'd73;  #10 
a = 8'd58; b = 8'd74;  #10 
a = 8'd58; b = 8'd75;  #10 
a = 8'd58; b = 8'd76;  #10 
a = 8'd58; b = 8'd77;  #10 
a = 8'd58; b = 8'd78;  #10 
a = 8'd58; b = 8'd79;  #10 
a = 8'd58; b = 8'd80;  #10 
a = 8'd58; b = 8'd81;  #10 
a = 8'd58; b = 8'd82;  #10 
a = 8'd58; b = 8'd83;  #10 
a = 8'd58; b = 8'd84;  #10 
a = 8'd58; b = 8'd85;  #10 
a = 8'd58; b = 8'd86;  #10 
a = 8'd58; b = 8'd87;  #10 
a = 8'd58; b = 8'd88;  #10 
a = 8'd58; b = 8'd89;  #10 
a = 8'd58; b = 8'd90;  #10 
a = 8'd58; b = 8'd91;  #10 
a = 8'd58; b = 8'd92;  #10 
a = 8'd58; b = 8'd93;  #10 
a = 8'd58; b = 8'd94;  #10 
a = 8'd58; b = 8'd95;  #10 
a = 8'd58; b = 8'd96;  #10 
a = 8'd58; b = 8'd97;  #10 
a = 8'd58; b = 8'd98;  #10 
a = 8'd58; b = 8'd99;  #10 
a = 8'd58; b = 8'd100;  #10 
a = 8'd58; b = 8'd101;  #10 
a = 8'd58; b = 8'd102;  #10 
a = 8'd58; b = 8'd103;  #10 
a = 8'd58; b = 8'd104;  #10 
a = 8'd58; b = 8'd105;  #10 
a = 8'd58; b = 8'd106;  #10 
a = 8'd58; b = 8'd107;  #10 
a = 8'd58; b = 8'd108;  #10 
a = 8'd58; b = 8'd109;  #10 
a = 8'd58; b = 8'd110;  #10 
a = 8'd58; b = 8'd111;  #10 
a = 8'd58; b = 8'd112;  #10 
a = 8'd58; b = 8'd113;  #10 
a = 8'd58; b = 8'd114;  #10 
a = 8'd58; b = 8'd115;  #10 
a = 8'd58; b = 8'd116;  #10 
a = 8'd58; b = 8'd117;  #10 
a = 8'd58; b = 8'd118;  #10 
a = 8'd58; b = 8'd119;  #10 
a = 8'd58; b = 8'd120;  #10 
a = 8'd58; b = 8'd121;  #10 
a = 8'd58; b = 8'd122;  #10 
a = 8'd58; b = 8'd123;  #10 
a = 8'd58; b = 8'd124;  #10 
a = 8'd58; b = 8'd125;  #10 
a = 8'd58; b = 8'd126;  #10 
a = 8'd58; b = 8'd127;  #10 
a = 8'd58; b = 8'd128;  #10 
a = 8'd58; b = 8'd129;  #10 
a = 8'd58; b = 8'd130;  #10 
a = 8'd58; b = 8'd131;  #10 
a = 8'd58; b = 8'd132;  #10 
a = 8'd58; b = 8'd133;  #10 
a = 8'd58; b = 8'd134;  #10 
a = 8'd58; b = 8'd135;  #10 
a = 8'd58; b = 8'd136;  #10 
a = 8'd58; b = 8'd137;  #10 
a = 8'd58; b = 8'd138;  #10 
a = 8'd58; b = 8'd139;  #10 
a = 8'd58; b = 8'd140;  #10 
a = 8'd58; b = 8'd141;  #10 
a = 8'd58; b = 8'd142;  #10 
a = 8'd58; b = 8'd143;  #10 
a = 8'd58; b = 8'd144;  #10 
a = 8'd58; b = 8'd145;  #10 
a = 8'd58; b = 8'd146;  #10 
a = 8'd58; b = 8'd147;  #10 
a = 8'd58; b = 8'd148;  #10 
a = 8'd58; b = 8'd149;  #10 
a = 8'd58; b = 8'd150;  #10 
a = 8'd58; b = 8'd151;  #10 
a = 8'd58; b = 8'd152;  #10 
a = 8'd58; b = 8'd153;  #10 
a = 8'd58; b = 8'd154;  #10 
a = 8'd58; b = 8'd155;  #10 
a = 8'd58; b = 8'd156;  #10 
a = 8'd58; b = 8'd157;  #10 
a = 8'd58; b = 8'd158;  #10 
a = 8'd58; b = 8'd159;  #10 
a = 8'd58; b = 8'd160;  #10 
a = 8'd58; b = 8'd161;  #10 
a = 8'd58; b = 8'd162;  #10 
a = 8'd58; b = 8'd163;  #10 
a = 8'd58; b = 8'd164;  #10 
a = 8'd58; b = 8'd165;  #10 
a = 8'd58; b = 8'd166;  #10 
a = 8'd58; b = 8'd167;  #10 
a = 8'd58; b = 8'd168;  #10 
a = 8'd58; b = 8'd169;  #10 
a = 8'd58; b = 8'd170;  #10 
a = 8'd58; b = 8'd171;  #10 
a = 8'd58; b = 8'd172;  #10 
a = 8'd58; b = 8'd173;  #10 
a = 8'd58; b = 8'd174;  #10 
a = 8'd58; b = 8'd175;  #10 
a = 8'd58; b = 8'd176;  #10 
a = 8'd58; b = 8'd177;  #10 
a = 8'd58; b = 8'd178;  #10 
a = 8'd58; b = 8'd179;  #10 
a = 8'd58; b = 8'd180;  #10 
a = 8'd58; b = 8'd181;  #10 
a = 8'd58; b = 8'd182;  #10 
a = 8'd58; b = 8'd183;  #10 
a = 8'd58; b = 8'd184;  #10 
a = 8'd58; b = 8'd185;  #10 
a = 8'd58; b = 8'd186;  #10 
a = 8'd58; b = 8'd187;  #10 
a = 8'd58; b = 8'd188;  #10 
a = 8'd58; b = 8'd189;  #10 
a = 8'd58; b = 8'd190;  #10 
a = 8'd58; b = 8'd191;  #10 
a = 8'd58; b = 8'd192;  #10 
a = 8'd58; b = 8'd193;  #10 
a = 8'd58; b = 8'd194;  #10 
a = 8'd58; b = 8'd195;  #10 
a = 8'd58; b = 8'd196;  #10 
a = 8'd58; b = 8'd197;  #10 
a = 8'd58; b = 8'd198;  #10 
a = 8'd58; b = 8'd199;  #10 
a = 8'd58; b = 8'd200;  #10 
a = 8'd58; b = 8'd201;  #10 
a = 8'd58; b = 8'd202;  #10 
a = 8'd58; b = 8'd203;  #10 
a = 8'd58; b = 8'd204;  #10 
a = 8'd58; b = 8'd205;  #10 
a = 8'd58; b = 8'd206;  #10 
a = 8'd58; b = 8'd207;  #10 
a = 8'd58; b = 8'd208;  #10 
a = 8'd58; b = 8'd209;  #10 
a = 8'd58; b = 8'd210;  #10 
a = 8'd58; b = 8'd211;  #10 
a = 8'd58; b = 8'd212;  #10 
a = 8'd58; b = 8'd213;  #10 
a = 8'd58; b = 8'd214;  #10 
a = 8'd58; b = 8'd215;  #10 
a = 8'd58; b = 8'd216;  #10 
a = 8'd58; b = 8'd217;  #10 
a = 8'd58; b = 8'd218;  #10 
a = 8'd58; b = 8'd219;  #10 
a = 8'd58; b = 8'd220;  #10 
a = 8'd58; b = 8'd221;  #10 
a = 8'd58; b = 8'd222;  #10 
a = 8'd58; b = 8'd223;  #10 
a = 8'd58; b = 8'd224;  #10 
a = 8'd58; b = 8'd225;  #10 
a = 8'd58; b = 8'd226;  #10 
a = 8'd58; b = 8'd227;  #10 
a = 8'd58; b = 8'd228;  #10 
a = 8'd58; b = 8'd229;  #10 
a = 8'd58; b = 8'd230;  #10 
a = 8'd58; b = 8'd231;  #10 
a = 8'd58; b = 8'd232;  #10 
a = 8'd58; b = 8'd233;  #10 
a = 8'd58; b = 8'd234;  #10 
a = 8'd58; b = 8'd235;  #10 
a = 8'd58; b = 8'd236;  #10 
a = 8'd58; b = 8'd237;  #10 
a = 8'd58; b = 8'd238;  #10 
a = 8'd58; b = 8'd239;  #10 
a = 8'd58; b = 8'd240;  #10 
a = 8'd58; b = 8'd241;  #10 
a = 8'd58; b = 8'd242;  #10 
a = 8'd58; b = 8'd243;  #10 
a = 8'd58; b = 8'd244;  #10 
a = 8'd58; b = 8'd245;  #10 
a = 8'd58; b = 8'd246;  #10 
a = 8'd58; b = 8'd247;  #10 
a = 8'd58; b = 8'd248;  #10 
a = 8'd58; b = 8'd249;  #10 
a = 8'd58; b = 8'd250;  #10 
a = 8'd58; b = 8'd251;  #10 
a = 8'd58; b = 8'd252;  #10 
a = 8'd58; b = 8'd253;  #10 
a = 8'd58; b = 8'd254;  #10 
a = 8'd58; b = 8'd255;  #10 
a = 8'd59; b = 8'd0;  #10 
a = 8'd59; b = 8'd1;  #10 
a = 8'd59; b = 8'd2;  #10 
a = 8'd59; b = 8'd3;  #10 
a = 8'd59; b = 8'd4;  #10 
a = 8'd59; b = 8'd5;  #10 
a = 8'd59; b = 8'd6;  #10 
a = 8'd59; b = 8'd7;  #10 
a = 8'd59; b = 8'd8;  #10 
a = 8'd59; b = 8'd9;  #10 
a = 8'd59; b = 8'd10;  #10 
a = 8'd59; b = 8'd11;  #10 
a = 8'd59; b = 8'd12;  #10 
a = 8'd59; b = 8'd13;  #10 
a = 8'd59; b = 8'd14;  #10 
a = 8'd59; b = 8'd15;  #10 
a = 8'd59; b = 8'd16;  #10 
a = 8'd59; b = 8'd17;  #10 
a = 8'd59; b = 8'd18;  #10 
a = 8'd59; b = 8'd19;  #10 
a = 8'd59; b = 8'd20;  #10 
a = 8'd59; b = 8'd21;  #10 
a = 8'd59; b = 8'd22;  #10 
a = 8'd59; b = 8'd23;  #10 
a = 8'd59; b = 8'd24;  #10 
a = 8'd59; b = 8'd25;  #10 
a = 8'd59; b = 8'd26;  #10 
a = 8'd59; b = 8'd27;  #10 
a = 8'd59; b = 8'd28;  #10 
a = 8'd59; b = 8'd29;  #10 
a = 8'd59; b = 8'd30;  #10 
a = 8'd59; b = 8'd31;  #10 
a = 8'd59; b = 8'd32;  #10 
a = 8'd59; b = 8'd33;  #10 
a = 8'd59; b = 8'd34;  #10 
a = 8'd59; b = 8'd35;  #10 
a = 8'd59; b = 8'd36;  #10 
a = 8'd59; b = 8'd37;  #10 
a = 8'd59; b = 8'd38;  #10 
a = 8'd59; b = 8'd39;  #10 
a = 8'd59; b = 8'd40;  #10 
a = 8'd59; b = 8'd41;  #10 
a = 8'd59; b = 8'd42;  #10 
a = 8'd59; b = 8'd43;  #10 
a = 8'd59; b = 8'd44;  #10 
a = 8'd59; b = 8'd45;  #10 
a = 8'd59; b = 8'd46;  #10 
a = 8'd59; b = 8'd47;  #10 
a = 8'd59; b = 8'd48;  #10 
a = 8'd59; b = 8'd49;  #10 
a = 8'd59; b = 8'd50;  #10 
a = 8'd59; b = 8'd51;  #10 
a = 8'd59; b = 8'd52;  #10 
a = 8'd59; b = 8'd53;  #10 
a = 8'd59; b = 8'd54;  #10 
a = 8'd59; b = 8'd55;  #10 
a = 8'd59; b = 8'd56;  #10 
a = 8'd59; b = 8'd57;  #10 
a = 8'd59; b = 8'd58;  #10 
a = 8'd59; b = 8'd59;  #10 
a = 8'd59; b = 8'd60;  #10 
a = 8'd59; b = 8'd61;  #10 
a = 8'd59; b = 8'd62;  #10 
a = 8'd59; b = 8'd63;  #10 
a = 8'd59; b = 8'd64;  #10 
a = 8'd59; b = 8'd65;  #10 
a = 8'd59; b = 8'd66;  #10 
a = 8'd59; b = 8'd67;  #10 
a = 8'd59; b = 8'd68;  #10 
a = 8'd59; b = 8'd69;  #10 
a = 8'd59; b = 8'd70;  #10 
a = 8'd59; b = 8'd71;  #10 
a = 8'd59; b = 8'd72;  #10 
a = 8'd59; b = 8'd73;  #10 
a = 8'd59; b = 8'd74;  #10 
a = 8'd59; b = 8'd75;  #10 
a = 8'd59; b = 8'd76;  #10 
a = 8'd59; b = 8'd77;  #10 
a = 8'd59; b = 8'd78;  #10 
a = 8'd59; b = 8'd79;  #10 
a = 8'd59; b = 8'd80;  #10 
a = 8'd59; b = 8'd81;  #10 
a = 8'd59; b = 8'd82;  #10 
a = 8'd59; b = 8'd83;  #10 
a = 8'd59; b = 8'd84;  #10 
a = 8'd59; b = 8'd85;  #10 
a = 8'd59; b = 8'd86;  #10 
a = 8'd59; b = 8'd87;  #10 
a = 8'd59; b = 8'd88;  #10 
a = 8'd59; b = 8'd89;  #10 
a = 8'd59; b = 8'd90;  #10 
a = 8'd59; b = 8'd91;  #10 
a = 8'd59; b = 8'd92;  #10 
a = 8'd59; b = 8'd93;  #10 
a = 8'd59; b = 8'd94;  #10 
a = 8'd59; b = 8'd95;  #10 
a = 8'd59; b = 8'd96;  #10 
a = 8'd59; b = 8'd97;  #10 
a = 8'd59; b = 8'd98;  #10 
a = 8'd59; b = 8'd99;  #10 
a = 8'd59; b = 8'd100;  #10 
a = 8'd59; b = 8'd101;  #10 
a = 8'd59; b = 8'd102;  #10 
a = 8'd59; b = 8'd103;  #10 
a = 8'd59; b = 8'd104;  #10 
a = 8'd59; b = 8'd105;  #10 
a = 8'd59; b = 8'd106;  #10 
a = 8'd59; b = 8'd107;  #10 
a = 8'd59; b = 8'd108;  #10 
a = 8'd59; b = 8'd109;  #10 
a = 8'd59; b = 8'd110;  #10 
a = 8'd59; b = 8'd111;  #10 
a = 8'd59; b = 8'd112;  #10 
a = 8'd59; b = 8'd113;  #10 
a = 8'd59; b = 8'd114;  #10 
a = 8'd59; b = 8'd115;  #10 
a = 8'd59; b = 8'd116;  #10 
a = 8'd59; b = 8'd117;  #10 
a = 8'd59; b = 8'd118;  #10 
a = 8'd59; b = 8'd119;  #10 
a = 8'd59; b = 8'd120;  #10 
a = 8'd59; b = 8'd121;  #10 
a = 8'd59; b = 8'd122;  #10 
a = 8'd59; b = 8'd123;  #10 
a = 8'd59; b = 8'd124;  #10 
a = 8'd59; b = 8'd125;  #10 
a = 8'd59; b = 8'd126;  #10 
a = 8'd59; b = 8'd127;  #10 
a = 8'd59; b = 8'd128;  #10 
a = 8'd59; b = 8'd129;  #10 
a = 8'd59; b = 8'd130;  #10 
a = 8'd59; b = 8'd131;  #10 
a = 8'd59; b = 8'd132;  #10 
a = 8'd59; b = 8'd133;  #10 
a = 8'd59; b = 8'd134;  #10 
a = 8'd59; b = 8'd135;  #10 
a = 8'd59; b = 8'd136;  #10 
a = 8'd59; b = 8'd137;  #10 
a = 8'd59; b = 8'd138;  #10 
a = 8'd59; b = 8'd139;  #10 
a = 8'd59; b = 8'd140;  #10 
a = 8'd59; b = 8'd141;  #10 
a = 8'd59; b = 8'd142;  #10 
a = 8'd59; b = 8'd143;  #10 
a = 8'd59; b = 8'd144;  #10 
a = 8'd59; b = 8'd145;  #10 
a = 8'd59; b = 8'd146;  #10 
a = 8'd59; b = 8'd147;  #10 
a = 8'd59; b = 8'd148;  #10 
a = 8'd59; b = 8'd149;  #10 
a = 8'd59; b = 8'd150;  #10 
a = 8'd59; b = 8'd151;  #10 
a = 8'd59; b = 8'd152;  #10 
a = 8'd59; b = 8'd153;  #10 
a = 8'd59; b = 8'd154;  #10 
a = 8'd59; b = 8'd155;  #10 
a = 8'd59; b = 8'd156;  #10 
a = 8'd59; b = 8'd157;  #10 
a = 8'd59; b = 8'd158;  #10 
a = 8'd59; b = 8'd159;  #10 
a = 8'd59; b = 8'd160;  #10 
a = 8'd59; b = 8'd161;  #10 
a = 8'd59; b = 8'd162;  #10 
a = 8'd59; b = 8'd163;  #10 
a = 8'd59; b = 8'd164;  #10 
a = 8'd59; b = 8'd165;  #10 
a = 8'd59; b = 8'd166;  #10 
a = 8'd59; b = 8'd167;  #10 
a = 8'd59; b = 8'd168;  #10 
a = 8'd59; b = 8'd169;  #10 
a = 8'd59; b = 8'd170;  #10 
a = 8'd59; b = 8'd171;  #10 
a = 8'd59; b = 8'd172;  #10 
a = 8'd59; b = 8'd173;  #10 
a = 8'd59; b = 8'd174;  #10 
a = 8'd59; b = 8'd175;  #10 
a = 8'd59; b = 8'd176;  #10 
a = 8'd59; b = 8'd177;  #10 
a = 8'd59; b = 8'd178;  #10 
a = 8'd59; b = 8'd179;  #10 
a = 8'd59; b = 8'd180;  #10 
a = 8'd59; b = 8'd181;  #10 
a = 8'd59; b = 8'd182;  #10 
a = 8'd59; b = 8'd183;  #10 
a = 8'd59; b = 8'd184;  #10 
a = 8'd59; b = 8'd185;  #10 
a = 8'd59; b = 8'd186;  #10 
a = 8'd59; b = 8'd187;  #10 
a = 8'd59; b = 8'd188;  #10 
a = 8'd59; b = 8'd189;  #10 
a = 8'd59; b = 8'd190;  #10 
a = 8'd59; b = 8'd191;  #10 
a = 8'd59; b = 8'd192;  #10 
a = 8'd59; b = 8'd193;  #10 
a = 8'd59; b = 8'd194;  #10 
a = 8'd59; b = 8'd195;  #10 
a = 8'd59; b = 8'd196;  #10 
a = 8'd59; b = 8'd197;  #10 
a = 8'd59; b = 8'd198;  #10 
a = 8'd59; b = 8'd199;  #10 
a = 8'd59; b = 8'd200;  #10 
a = 8'd59; b = 8'd201;  #10 
a = 8'd59; b = 8'd202;  #10 
a = 8'd59; b = 8'd203;  #10 
a = 8'd59; b = 8'd204;  #10 
a = 8'd59; b = 8'd205;  #10 
a = 8'd59; b = 8'd206;  #10 
a = 8'd59; b = 8'd207;  #10 
a = 8'd59; b = 8'd208;  #10 
a = 8'd59; b = 8'd209;  #10 
a = 8'd59; b = 8'd210;  #10 
a = 8'd59; b = 8'd211;  #10 
a = 8'd59; b = 8'd212;  #10 
a = 8'd59; b = 8'd213;  #10 
a = 8'd59; b = 8'd214;  #10 
a = 8'd59; b = 8'd215;  #10 
a = 8'd59; b = 8'd216;  #10 
a = 8'd59; b = 8'd217;  #10 
a = 8'd59; b = 8'd218;  #10 
a = 8'd59; b = 8'd219;  #10 
a = 8'd59; b = 8'd220;  #10 
a = 8'd59; b = 8'd221;  #10 
a = 8'd59; b = 8'd222;  #10 
a = 8'd59; b = 8'd223;  #10 
a = 8'd59; b = 8'd224;  #10 
a = 8'd59; b = 8'd225;  #10 
a = 8'd59; b = 8'd226;  #10 
a = 8'd59; b = 8'd227;  #10 
a = 8'd59; b = 8'd228;  #10 
a = 8'd59; b = 8'd229;  #10 
a = 8'd59; b = 8'd230;  #10 
a = 8'd59; b = 8'd231;  #10 
a = 8'd59; b = 8'd232;  #10 
a = 8'd59; b = 8'd233;  #10 
a = 8'd59; b = 8'd234;  #10 
a = 8'd59; b = 8'd235;  #10 
a = 8'd59; b = 8'd236;  #10 
a = 8'd59; b = 8'd237;  #10 
a = 8'd59; b = 8'd238;  #10 
a = 8'd59; b = 8'd239;  #10 
a = 8'd59; b = 8'd240;  #10 
a = 8'd59; b = 8'd241;  #10 
a = 8'd59; b = 8'd242;  #10 
a = 8'd59; b = 8'd243;  #10 
a = 8'd59; b = 8'd244;  #10 
a = 8'd59; b = 8'd245;  #10 
a = 8'd59; b = 8'd246;  #10 
a = 8'd59; b = 8'd247;  #10 
a = 8'd59; b = 8'd248;  #10 
a = 8'd59; b = 8'd249;  #10 
a = 8'd59; b = 8'd250;  #10 
a = 8'd59; b = 8'd251;  #10 
a = 8'd59; b = 8'd252;  #10 
a = 8'd59; b = 8'd253;  #10 
a = 8'd59; b = 8'd254;  #10 
a = 8'd59; b = 8'd255;  #10 
a = 8'd60; b = 8'd0;  #10 
a = 8'd60; b = 8'd1;  #10 
a = 8'd60; b = 8'd2;  #10 
a = 8'd60; b = 8'd3;  #10 
a = 8'd60; b = 8'd4;  #10 
a = 8'd60; b = 8'd5;  #10 
a = 8'd60; b = 8'd6;  #10 
a = 8'd60; b = 8'd7;  #10 
a = 8'd60; b = 8'd8;  #10 
a = 8'd60; b = 8'd9;  #10 
a = 8'd60; b = 8'd10;  #10 
a = 8'd60; b = 8'd11;  #10 
a = 8'd60; b = 8'd12;  #10 
a = 8'd60; b = 8'd13;  #10 
a = 8'd60; b = 8'd14;  #10 
a = 8'd60; b = 8'd15;  #10 
a = 8'd60; b = 8'd16;  #10 
a = 8'd60; b = 8'd17;  #10 
a = 8'd60; b = 8'd18;  #10 
a = 8'd60; b = 8'd19;  #10 
a = 8'd60; b = 8'd20;  #10 
a = 8'd60; b = 8'd21;  #10 
a = 8'd60; b = 8'd22;  #10 
a = 8'd60; b = 8'd23;  #10 
a = 8'd60; b = 8'd24;  #10 
a = 8'd60; b = 8'd25;  #10 
a = 8'd60; b = 8'd26;  #10 
a = 8'd60; b = 8'd27;  #10 
a = 8'd60; b = 8'd28;  #10 
a = 8'd60; b = 8'd29;  #10 
a = 8'd60; b = 8'd30;  #10 
a = 8'd60; b = 8'd31;  #10 
a = 8'd60; b = 8'd32;  #10 
a = 8'd60; b = 8'd33;  #10 
a = 8'd60; b = 8'd34;  #10 
a = 8'd60; b = 8'd35;  #10 
a = 8'd60; b = 8'd36;  #10 
a = 8'd60; b = 8'd37;  #10 
a = 8'd60; b = 8'd38;  #10 
a = 8'd60; b = 8'd39;  #10 
a = 8'd60; b = 8'd40;  #10 
a = 8'd60; b = 8'd41;  #10 
a = 8'd60; b = 8'd42;  #10 
a = 8'd60; b = 8'd43;  #10 
a = 8'd60; b = 8'd44;  #10 
a = 8'd60; b = 8'd45;  #10 
a = 8'd60; b = 8'd46;  #10 
a = 8'd60; b = 8'd47;  #10 
a = 8'd60; b = 8'd48;  #10 
a = 8'd60; b = 8'd49;  #10 
a = 8'd60; b = 8'd50;  #10 
a = 8'd60; b = 8'd51;  #10 
a = 8'd60; b = 8'd52;  #10 
a = 8'd60; b = 8'd53;  #10 
a = 8'd60; b = 8'd54;  #10 
a = 8'd60; b = 8'd55;  #10 
a = 8'd60; b = 8'd56;  #10 
a = 8'd60; b = 8'd57;  #10 
a = 8'd60; b = 8'd58;  #10 
a = 8'd60; b = 8'd59;  #10 
a = 8'd60; b = 8'd60;  #10 
a = 8'd60; b = 8'd61;  #10 
a = 8'd60; b = 8'd62;  #10 
a = 8'd60; b = 8'd63;  #10 
a = 8'd60; b = 8'd64;  #10 
a = 8'd60; b = 8'd65;  #10 
a = 8'd60; b = 8'd66;  #10 
a = 8'd60; b = 8'd67;  #10 
a = 8'd60; b = 8'd68;  #10 
a = 8'd60; b = 8'd69;  #10 
a = 8'd60; b = 8'd70;  #10 
a = 8'd60; b = 8'd71;  #10 
a = 8'd60; b = 8'd72;  #10 
a = 8'd60; b = 8'd73;  #10 
a = 8'd60; b = 8'd74;  #10 
a = 8'd60; b = 8'd75;  #10 
a = 8'd60; b = 8'd76;  #10 
a = 8'd60; b = 8'd77;  #10 
a = 8'd60; b = 8'd78;  #10 
a = 8'd60; b = 8'd79;  #10 
a = 8'd60; b = 8'd80;  #10 
a = 8'd60; b = 8'd81;  #10 
a = 8'd60; b = 8'd82;  #10 
a = 8'd60; b = 8'd83;  #10 
a = 8'd60; b = 8'd84;  #10 
a = 8'd60; b = 8'd85;  #10 
a = 8'd60; b = 8'd86;  #10 
a = 8'd60; b = 8'd87;  #10 
a = 8'd60; b = 8'd88;  #10 
a = 8'd60; b = 8'd89;  #10 
a = 8'd60; b = 8'd90;  #10 
a = 8'd60; b = 8'd91;  #10 
a = 8'd60; b = 8'd92;  #10 
a = 8'd60; b = 8'd93;  #10 
a = 8'd60; b = 8'd94;  #10 
a = 8'd60; b = 8'd95;  #10 
a = 8'd60; b = 8'd96;  #10 
a = 8'd60; b = 8'd97;  #10 
a = 8'd60; b = 8'd98;  #10 
a = 8'd60; b = 8'd99;  #10 
a = 8'd60; b = 8'd100;  #10 
a = 8'd60; b = 8'd101;  #10 
a = 8'd60; b = 8'd102;  #10 
a = 8'd60; b = 8'd103;  #10 
a = 8'd60; b = 8'd104;  #10 
a = 8'd60; b = 8'd105;  #10 
a = 8'd60; b = 8'd106;  #10 
a = 8'd60; b = 8'd107;  #10 
a = 8'd60; b = 8'd108;  #10 
a = 8'd60; b = 8'd109;  #10 
a = 8'd60; b = 8'd110;  #10 
a = 8'd60; b = 8'd111;  #10 
a = 8'd60; b = 8'd112;  #10 
a = 8'd60; b = 8'd113;  #10 
a = 8'd60; b = 8'd114;  #10 
a = 8'd60; b = 8'd115;  #10 
a = 8'd60; b = 8'd116;  #10 
a = 8'd60; b = 8'd117;  #10 
a = 8'd60; b = 8'd118;  #10 
a = 8'd60; b = 8'd119;  #10 
a = 8'd60; b = 8'd120;  #10 
a = 8'd60; b = 8'd121;  #10 
a = 8'd60; b = 8'd122;  #10 
a = 8'd60; b = 8'd123;  #10 
a = 8'd60; b = 8'd124;  #10 
a = 8'd60; b = 8'd125;  #10 
a = 8'd60; b = 8'd126;  #10 
a = 8'd60; b = 8'd127;  #10 
a = 8'd60; b = 8'd128;  #10 
a = 8'd60; b = 8'd129;  #10 
a = 8'd60; b = 8'd130;  #10 
a = 8'd60; b = 8'd131;  #10 
a = 8'd60; b = 8'd132;  #10 
a = 8'd60; b = 8'd133;  #10 
a = 8'd60; b = 8'd134;  #10 
a = 8'd60; b = 8'd135;  #10 
a = 8'd60; b = 8'd136;  #10 
a = 8'd60; b = 8'd137;  #10 
a = 8'd60; b = 8'd138;  #10 
a = 8'd60; b = 8'd139;  #10 
a = 8'd60; b = 8'd140;  #10 
a = 8'd60; b = 8'd141;  #10 
a = 8'd60; b = 8'd142;  #10 
a = 8'd60; b = 8'd143;  #10 
a = 8'd60; b = 8'd144;  #10 
a = 8'd60; b = 8'd145;  #10 
a = 8'd60; b = 8'd146;  #10 
a = 8'd60; b = 8'd147;  #10 
a = 8'd60; b = 8'd148;  #10 
a = 8'd60; b = 8'd149;  #10 
a = 8'd60; b = 8'd150;  #10 
a = 8'd60; b = 8'd151;  #10 
a = 8'd60; b = 8'd152;  #10 
a = 8'd60; b = 8'd153;  #10 
a = 8'd60; b = 8'd154;  #10 
a = 8'd60; b = 8'd155;  #10 
a = 8'd60; b = 8'd156;  #10 
a = 8'd60; b = 8'd157;  #10 
a = 8'd60; b = 8'd158;  #10 
a = 8'd60; b = 8'd159;  #10 
a = 8'd60; b = 8'd160;  #10 
a = 8'd60; b = 8'd161;  #10 
a = 8'd60; b = 8'd162;  #10 
a = 8'd60; b = 8'd163;  #10 
a = 8'd60; b = 8'd164;  #10 
a = 8'd60; b = 8'd165;  #10 
a = 8'd60; b = 8'd166;  #10 
a = 8'd60; b = 8'd167;  #10 
a = 8'd60; b = 8'd168;  #10 
a = 8'd60; b = 8'd169;  #10 
a = 8'd60; b = 8'd170;  #10 
a = 8'd60; b = 8'd171;  #10 
a = 8'd60; b = 8'd172;  #10 
a = 8'd60; b = 8'd173;  #10 
a = 8'd60; b = 8'd174;  #10 
a = 8'd60; b = 8'd175;  #10 
a = 8'd60; b = 8'd176;  #10 
a = 8'd60; b = 8'd177;  #10 
a = 8'd60; b = 8'd178;  #10 
a = 8'd60; b = 8'd179;  #10 
a = 8'd60; b = 8'd180;  #10 
a = 8'd60; b = 8'd181;  #10 
a = 8'd60; b = 8'd182;  #10 
a = 8'd60; b = 8'd183;  #10 
a = 8'd60; b = 8'd184;  #10 
a = 8'd60; b = 8'd185;  #10 
a = 8'd60; b = 8'd186;  #10 
a = 8'd60; b = 8'd187;  #10 
a = 8'd60; b = 8'd188;  #10 
a = 8'd60; b = 8'd189;  #10 
a = 8'd60; b = 8'd190;  #10 
a = 8'd60; b = 8'd191;  #10 
a = 8'd60; b = 8'd192;  #10 
a = 8'd60; b = 8'd193;  #10 
a = 8'd60; b = 8'd194;  #10 
a = 8'd60; b = 8'd195;  #10 
a = 8'd60; b = 8'd196;  #10 
a = 8'd60; b = 8'd197;  #10 
a = 8'd60; b = 8'd198;  #10 
a = 8'd60; b = 8'd199;  #10 
a = 8'd60; b = 8'd200;  #10 
a = 8'd60; b = 8'd201;  #10 
a = 8'd60; b = 8'd202;  #10 
a = 8'd60; b = 8'd203;  #10 
a = 8'd60; b = 8'd204;  #10 
a = 8'd60; b = 8'd205;  #10 
a = 8'd60; b = 8'd206;  #10 
a = 8'd60; b = 8'd207;  #10 
a = 8'd60; b = 8'd208;  #10 
a = 8'd60; b = 8'd209;  #10 
a = 8'd60; b = 8'd210;  #10 
a = 8'd60; b = 8'd211;  #10 
a = 8'd60; b = 8'd212;  #10 
a = 8'd60; b = 8'd213;  #10 
a = 8'd60; b = 8'd214;  #10 
a = 8'd60; b = 8'd215;  #10 
a = 8'd60; b = 8'd216;  #10 
a = 8'd60; b = 8'd217;  #10 
a = 8'd60; b = 8'd218;  #10 
a = 8'd60; b = 8'd219;  #10 
a = 8'd60; b = 8'd220;  #10 
a = 8'd60; b = 8'd221;  #10 
a = 8'd60; b = 8'd222;  #10 
a = 8'd60; b = 8'd223;  #10 
a = 8'd60; b = 8'd224;  #10 
a = 8'd60; b = 8'd225;  #10 
a = 8'd60; b = 8'd226;  #10 
a = 8'd60; b = 8'd227;  #10 
a = 8'd60; b = 8'd228;  #10 
a = 8'd60; b = 8'd229;  #10 
a = 8'd60; b = 8'd230;  #10 
a = 8'd60; b = 8'd231;  #10 
a = 8'd60; b = 8'd232;  #10 
a = 8'd60; b = 8'd233;  #10 
a = 8'd60; b = 8'd234;  #10 
a = 8'd60; b = 8'd235;  #10 
a = 8'd60; b = 8'd236;  #10 
a = 8'd60; b = 8'd237;  #10 
a = 8'd60; b = 8'd238;  #10 
a = 8'd60; b = 8'd239;  #10 
a = 8'd60; b = 8'd240;  #10 
a = 8'd60; b = 8'd241;  #10 
a = 8'd60; b = 8'd242;  #10 
a = 8'd60; b = 8'd243;  #10 
a = 8'd60; b = 8'd244;  #10 
a = 8'd60; b = 8'd245;  #10 
a = 8'd60; b = 8'd246;  #10 
a = 8'd60; b = 8'd247;  #10 
a = 8'd60; b = 8'd248;  #10 
a = 8'd60; b = 8'd249;  #10 
a = 8'd60; b = 8'd250;  #10 
a = 8'd60; b = 8'd251;  #10 
a = 8'd60; b = 8'd252;  #10 
a = 8'd60; b = 8'd253;  #10 
a = 8'd60; b = 8'd254;  #10 
a = 8'd60; b = 8'd255;  #10 
a = 8'd61; b = 8'd0;  #10 
a = 8'd61; b = 8'd1;  #10 
a = 8'd61; b = 8'd2;  #10 
a = 8'd61; b = 8'd3;  #10 
a = 8'd61; b = 8'd4;  #10 
a = 8'd61; b = 8'd5;  #10 
a = 8'd61; b = 8'd6;  #10 
a = 8'd61; b = 8'd7;  #10 
a = 8'd61; b = 8'd8;  #10 
a = 8'd61; b = 8'd9;  #10 
a = 8'd61; b = 8'd10;  #10 
a = 8'd61; b = 8'd11;  #10 
a = 8'd61; b = 8'd12;  #10 
a = 8'd61; b = 8'd13;  #10 
a = 8'd61; b = 8'd14;  #10 
a = 8'd61; b = 8'd15;  #10 
a = 8'd61; b = 8'd16;  #10 
a = 8'd61; b = 8'd17;  #10 
a = 8'd61; b = 8'd18;  #10 
a = 8'd61; b = 8'd19;  #10 
a = 8'd61; b = 8'd20;  #10 
a = 8'd61; b = 8'd21;  #10 
a = 8'd61; b = 8'd22;  #10 
a = 8'd61; b = 8'd23;  #10 
a = 8'd61; b = 8'd24;  #10 
a = 8'd61; b = 8'd25;  #10 
a = 8'd61; b = 8'd26;  #10 
a = 8'd61; b = 8'd27;  #10 
a = 8'd61; b = 8'd28;  #10 
a = 8'd61; b = 8'd29;  #10 
a = 8'd61; b = 8'd30;  #10 
a = 8'd61; b = 8'd31;  #10 
a = 8'd61; b = 8'd32;  #10 
a = 8'd61; b = 8'd33;  #10 
a = 8'd61; b = 8'd34;  #10 
a = 8'd61; b = 8'd35;  #10 
a = 8'd61; b = 8'd36;  #10 
a = 8'd61; b = 8'd37;  #10 
a = 8'd61; b = 8'd38;  #10 
a = 8'd61; b = 8'd39;  #10 
a = 8'd61; b = 8'd40;  #10 
a = 8'd61; b = 8'd41;  #10 
a = 8'd61; b = 8'd42;  #10 
a = 8'd61; b = 8'd43;  #10 
a = 8'd61; b = 8'd44;  #10 
a = 8'd61; b = 8'd45;  #10 
a = 8'd61; b = 8'd46;  #10 
a = 8'd61; b = 8'd47;  #10 
a = 8'd61; b = 8'd48;  #10 
a = 8'd61; b = 8'd49;  #10 
a = 8'd61; b = 8'd50;  #10 
a = 8'd61; b = 8'd51;  #10 
a = 8'd61; b = 8'd52;  #10 
a = 8'd61; b = 8'd53;  #10 
a = 8'd61; b = 8'd54;  #10 
a = 8'd61; b = 8'd55;  #10 
a = 8'd61; b = 8'd56;  #10 
a = 8'd61; b = 8'd57;  #10 
a = 8'd61; b = 8'd58;  #10 
a = 8'd61; b = 8'd59;  #10 
a = 8'd61; b = 8'd60;  #10 
a = 8'd61; b = 8'd61;  #10 
a = 8'd61; b = 8'd62;  #10 
a = 8'd61; b = 8'd63;  #10 
a = 8'd61; b = 8'd64;  #10 
a = 8'd61; b = 8'd65;  #10 
a = 8'd61; b = 8'd66;  #10 
a = 8'd61; b = 8'd67;  #10 
a = 8'd61; b = 8'd68;  #10 
a = 8'd61; b = 8'd69;  #10 
a = 8'd61; b = 8'd70;  #10 
a = 8'd61; b = 8'd71;  #10 
a = 8'd61; b = 8'd72;  #10 
a = 8'd61; b = 8'd73;  #10 
a = 8'd61; b = 8'd74;  #10 
a = 8'd61; b = 8'd75;  #10 
a = 8'd61; b = 8'd76;  #10 
a = 8'd61; b = 8'd77;  #10 
a = 8'd61; b = 8'd78;  #10 
a = 8'd61; b = 8'd79;  #10 
a = 8'd61; b = 8'd80;  #10 
a = 8'd61; b = 8'd81;  #10 
a = 8'd61; b = 8'd82;  #10 
a = 8'd61; b = 8'd83;  #10 
a = 8'd61; b = 8'd84;  #10 
a = 8'd61; b = 8'd85;  #10 
a = 8'd61; b = 8'd86;  #10 
a = 8'd61; b = 8'd87;  #10 
a = 8'd61; b = 8'd88;  #10 
a = 8'd61; b = 8'd89;  #10 
a = 8'd61; b = 8'd90;  #10 
a = 8'd61; b = 8'd91;  #10 
a = 8'd61; b = 8'd92;  #10 
a = 8'd61; b = 8'd93;  #10 
a = 8'd61; b = 8'd94;  #10 
a = 8'd61; b = 8'd95;  #10 
a = 8'd61; b = 8'd96;  #10 
a = 8'd61; b = 8'd97;  #10 
a = 8'd61; b = 8'd98;  #10 
a = 8'd61; b = 8'd99;  #10 
a = 8'd61; b = 8'd100;  #10 
a = 8'd61; b = 8'd101;  #10 
a = 8'd61; b = 8'd102;  #10 
a = 8'd61; b = 8'd103;  #10 
a = 8'd61; b = 8'd104;  #10 
a = 8'd61; b = 8'd105;  #10 
a = 8'd61; b = 8'd106;  #10 
a = 8'd61; b = 8'd107;  #10 
a = 8'd61; b = 8'd108;  #10 
a = 8'd61; b = 8'd109;  #10 
a = 8'd61; b = 8'd110;  #10 
a = 8'd61; b = 8'd111;  #10 
a = 8'd61; b = 8'd112;  #10 
a = 8'd61; b = 8'd113;  #10 
a = 8'd61; b = 8'd114;  #10 
a = 8'd61; b = 8'd115;  #10 
a = 8'd61; b = 8'd116;  #10 
a = 8'd61; b = 8'd117;  #10 
a = 8'd61; b = 8'd118;  #10 
a = 8'd61; b = 8'd119;  #10 
a = 8'd61; b = 8'd120;  #10 
a = 8'd61; b = 8'd121;  #10 
a = 8'd61; b = 8'd122;  #10 
a = 8'd61; b = 8'd123;  #10 
a = 8'd61; b = 8'd124;  #10 
a = 8'd61; b = 8'd125;  #10 
a = 8'd61; b = 8'd126;  #10 
a = 8'd61; b = 8'd127;  #10 
a = 8'd61; b = 8'd128;  #10 
a = 8'd61; b = 8'd129;  #10 
a = 8'd61; b = 8'd130;  #10 
a = 8'd61; b = 8'd131;  #10 
a = 8'd61; b = 8'd132;  #10 
a = 8'd61; b = 8'd133;  #10 
a = 8'd61; b = 8'd134;  #10 
a = 8'd61; b = 8'd135;  #10 
a = 8'd61; b = 8'd136;  #10 
a = 8'd61; b = 8'd137;  #10 
a = 8'd61; b = 8'd138;  #10 
a = 8'd61; b = 8'd139;  #10 
a = 8'd61; b = 8'd140;  #10 
a = 8'd61; b = 8'd141;  #10 
a = 8'd61; b = 8'd142;  #10 
a = 8'd61; b = 8'd143;  #10 
a = 8'd61; b = 8'd144;  #10 
a = 8'd61; b = 8'd145;  #10 
a = 8'd61; b = 8'd146;  #10 
a = 8'd61; b = 8'd147;  #10 
a = 8'd61; b = 8'd148;  #10 
a = 8'd61; b = 8'd149;  #10 
a = 8'd61; b = 8'd150;  #10 
a = 8'd61; b = 8'd151;  #10 
a = 8'd61; b = 8'd152;  #10 
a = 8'd61; b = 8'd153;  #10 
a = 8'd61; b = 8'd154;  #10 
a = 8'd61; b = 8'd155;  #10 
a = 8'd61; b = 8'd156;  #10 
a = 8'd61; b = 8'd157;  #10 
a = 8'd61; b = 8'd158;  #10 
a = 8'd61; b = 8'd159;  #10 
a = 8'd61; b = 8'd160;  #10 
a = 8'd61; b = 8'd161;  #10 
a = 8'd61; b = 8'd162;  #10 
a = 8'd61; b = 8'd163;  #10 
a = 8'd61; b = 8'd164;  #10 
a = 8'd61; b = 8'd165;  #10 
a = 8'd61; b = 8'd166;  #10 
a = 8'd61; b = 8'd167;  #10 
a = 8'd61; b = 8'd168;  #10 
a = 8'd61; b = 8'd169;  #10 
a = 8'd61; b = 8'd170;  #10 
a = 8'd61; b = 8'd171;  #10 
a = 8'd61; b = 8'd172;  #10 
a = 8'd61; b = 8'd173;  #10 
a = 8'd61; b = 8'd174;  #10 
a = 8'd61; b = 8'd175;  #10 
a = 8'd61; b = 8'd176;  #10 
a = 8'd61; b = 8'd177;  #10 
a = 8'd61; b = 8'd178;  #10 
a = 8'd61; b = 8'd179;  #10 
a = 8'd61; b = 8'd180;  #10 
a = 8'd61; b = 8'd181;  #10 
a = 8'd61; b = 8'd182;  #10 
a = 8'd61; b = 8'd183;  #10 
a = 8'd61; b = 8'd184;  #10 
a = 8'd61; b = 8'd185;  #10 
a = 8'd61; b = 8'd186;  #10 
a = 8'd61; b = 8'd187;  #10 
a = 8'd61; b = 8'd188;  #10 
a = 8'd61; b = 8'd189;  #10 
a = 8'd61; b = 8'd190;  #10 
a = 8'd61; b = 8'd191;  #10 
a = 8'd61; b = 8'd192;  #10 
a = 8'd61; b = 8'd193;  #10 
a = 8'd61; b = 8'd194;  #10 
a = 8'd61; b = 8'd195;  #10 
a = 8'd61; b = 8'd196;  #10 
a = 8'd61; b = 8'd197;  #10 
a = 8'd61; b = 8'd198;  #10 
a = 8'd61; b = 8'd199;  #10 
a = 8'd61; b = 8'd200;  #10 
a = 8'd61; b = 8'd201;  #10 
a = 8'd61; b = 8'd202;  #10 
a = 8'd61; b = 8'd203;  #10 
a = 8'd61; b = 8'd204;  #10 
a = 8'd61; b = 8'd205;  #10 
a = 8'd61; b = 8'd206;  #10 
a = 8'd61; b = 8'd207;  #10 
a = 8'd61; b = 8'd208;  #10 
a = 8'd61; b = 8'd209;  #10 
a = 8'd61; b = 8'd210;  #10 
a = 8'd61; b = 8'd211;  #10 
a = 8'd61; b = 8'd212;  #10 
a = 8'd61; b = 8'd213;  #10 
a = 8'd61; b = 8'd214;  #10 
a = 8'd61; b = 8'd215;  #10 
a = 8'd61; b = 8'd216;  #10 
a = 8'd61; b = 8'd217;  #10 
a = 8'd61; b = 8'd218;  #10 
a = 8'd61; b = 8'd219;  #10 
a = 8'd61; b = 8'd220;  #10 
a = 8'd61; b = 8'd221;  #10 
a = 8'd61; b = 8'd222;  #10 
a = 8'd61; b = 8'd223;  #10 
a = 8'd61; b = 8'd224;  #10 
a = 8'd61; b = 8'd225;  #10 
a = 8'd61; b = 8'd226;  #10 
a = 8'd61; b = 8'd227;  #10 
a = 8'd61; b = 8'd228;  #10 
a = 8'd61; b = 8'd229;  #10 
a = 8'd61; b = 8'd230;  #10 
a = 8'd61; b = 8'd231;  #10 
a = 8'd61; b = 8'd232;  #10 
a = 8'd61; b = 8'd233;  #10 
a = 8'd61; b = 8'd234;  #10 
a = 8'd61; b = 8'd235;  #10 
a = 8'd61; b = 8'd236;  #10 
a = 8'd61; b = 8'd237;  #10 
a = 8'd61; b = 8'd238;  #10 
a = 8'd61; b = 8'd239;  #10 
a = 8'd61; b = 8'd240;  #10 
a = 8'd61; b = 8'd241;  #10 
a = 8'd61; b = 8'd242;  #10 
a = 8'd61; b = 8'd243;  #10 
a = 8'd61; b = 8'd244;  #10 
a = 8'd61; b = 8'd245;  #10 
a = 8'd61; b = 8'd246;  #10 
a = 8'd61; b = 8'd247;  #10 
a = 8'd61; b = 8'd248;  #10 
a = 8'd61; b = 8'd249;  #10 
a = 8'd61; b = 8'd250;  #10 
a = 8'd61; b = 8'd251;  #10 
a = 8'd61; b = 8'd252;  #10 
a = 8'd61; b = 8'd253;  #10 
a = 8'd61; b = 8'd254;  #10 
a = 8'd61; b = 8'd255;  #10 
a = 8'd62; b = 8'd0;  #10 
a = 8'd62; b = 8'd1;  #10 
a = 8'd62; b = 8'd2;  #10 
a = 8'd62; b = 8'd3;  #10 
a = 8'd62; b = 8'd4;  #10 
a = 8'd62; b = 8'd5;  #10 
a = 8'd62; b = 8'd6;  #10 
a = 8'd62; b = 8'd7;  #10 
a = 8'd62; b = 8'd8;  #10 
a = 8'd62; b = 8'd9;  #10 
a = 8'd62; b = 8'd10;  #10 
a = 8'd62; b = 8'd11;  #10 
a = 8'd62; b = 8'd12;  #10 
a = 8'd62; b = 8'd13;  #10 
a = 8'd62; b = 8'd14;  #10 
a = 8'd62; b = 8'd15;  #10 
a = 8'd62; b = 8'd16;  #10 
a = 8'd62; b = 8'd17;  #10 
a = 8'd62; b = 8'd18;  #10 
a = 8'd62; b = 8'd19;  #10 
a = 8'd62; b = 8'd20;  #10 
a = 8'd62; b = 8'd21;  #10 
a = 8'd62; b = 8'd22;  #10 
a = 8'd62; b = 8'd23;  #10 
a = 8'd62; b = 8'd24;  #10 
a = 8'd62; b = 8'd25;  #10 
a = 8'd62; b = 8'd26;  #10 
a = 8'd62; b = 8'd27;  #10 
a = 8'd62; b = 8'd28;  #10 
a = 8'd62; b = 8'd29;  #10 
a = 8'd62; b = 8'd30;  #10 
a = 8'd62; b = 8'd31;  #10 
a = 8'd62; b = 8'd32;  #10 
a = 8'd62; b = 8'd33;  #10 
a = 8'd62; b = 8'd34;  #10 
a = 8'd62; b = 8'd35;  #10 
a = 8'd62; b = 8'd36;  #10 
a = 8'd62; b = 8'd37;  #10 
a = 8'd62; b = 8'd38;  #10 
a = 8'd62; b = 8'd39;  #10 
a = 8'd62; b = 8'd40;  #10 
a = 8'd62; b = 8'd41;  #10 
a = 8'd62; b = 8'd42;  #10 
a = 8'd62; b = 8'd43;  #10 
a = 8'd62; b = 8'd44;  #10 
a = 8'd62; b = 8'd45;  #10 
a = 8'd62; b = 8'd46;  #10 
a = 8'd62; b = 8'd47;  #10 
a = 8'd62; b = 8'd48;  #10 
a = 8'd62; b = 8'd49;  #10 
a = 8'd62; b = 8'd50;  #10 
a = 8'd62; b = 8'd51;  #10 
a = 8'd62; b = 8'd52;  #10 
a = 8'd62; b = 8'd53;  #10 
a = 8'd62; b = 8'd54;  #10 
a = 8'd62; b = 8'd55;  #10 
a = 8'd62; b = 8'd56;  #10 
a = 8'd62; b = 8'd57;  #10 
a = 8'd62; b = 8'd58;  #10 
a = 8'd62; b = 8'd59;  #10 
a = 8'd62; b = 8'd60;  #10 
a = 8'd62; b = 8'd61;  #10 
a = 8'd62; b = 8'd62;  #10 
a = 8'd62; b = 8'd63;  #10 
a = 8'd62; b = 8'd64;  #10 
a = 8'd62; b = 8'd65;  #10 
a = 8'd62; b = 8'd66;  #10 
a = 8'd62; b = 8'd67;  #10 
a = 8'd62; b = 8'd68;  #10 
a = 8'd62; b = 8'd69;  #10 
a = 8'd62; b = 8'd70;  #10 
a = 8'd62; b = 8'd71;  #10 
a = 8'd62; b = 8'd72;  #10 
a = 8'd62; b = 8'd73;  #10 
a = 8'd62; b = 8'd74;  #10 
a = 8'd62; b = 8'd75;  #10 
a = 8'd62; b = 8'd76;  #10 
a = 8'd62; b = 8'd77;  #10 
a = 8'd62; b = 8'd78;  #10 
a = 8'd62; b = 8'd79;  #10 
a = 8'd62; b = 8'd80;  #10 
a = 8'd62; b = 8'd81;  #10 
a = 8'd62; b = 8'd82;  #10 
a = 8'd62; b = 8'd83;  #10 
a = 8'd62; b = 8'd84;  #10 
a = 8'd62; b = 8'd85;  #10 
a = 8'd62; b = 8'd86;  #10 
a = 8'd62; b = 8'd87;  #10 
a = 8'd62; b = 8'd88;  #10 
a = 8'd62; b = 8'd89;  #10 
a = 8'd62; b = 8'd90;  #10 
a = 8'd62; b = 8'd91;  #10 
a = 8'd62; b = 8'd92;  #10 
a = 8'd62; b = 8'd93;  #10 
a = 8'd62; b = 8'd94;  #10 
a = 8'd62; b = 8'd95;  #10 
a = 8'd62; b = 8'd96;  #10 
a = 8'd62; b = 8'd97;  #10 
a = 8'd62; b = 8'd98;  #10 
a = 8'd62; b = 8'd99;  #10 
a = 8'd62; b = 8'd100;  #10 
a = 8'd62; b = 8'd101;  #10 
a = 8'd62; b = 8'd102;  #10 
a = 8'd62; b = 8'd103;  #10 
a = 8'd62; b = 8'd104;  #10 
a = 8'd62; b = 8'd105;  #10 
a = 8'd62; b = 8'd106;  #10 
a = 8'd62; b = 8'd107;  #10 
a = 8'd62; b = 8'd108;  #10 
a = 8'd62; b = 8'd109;  #10 
a = 8'd62; b = 8'd110;  #10 
a = 8'd62; b = 8'd111;  #10 
a = 8'd62; b = 8'd112;  #10 
a = 8'd62; b = 8'd113;  #10 
a = 8'd62; b = 8'd114;  #10 
a = 8'd62; b = 8'd115;  #10 
a = 8'd62; b = 8'd116;  #10 
a = 8'd62; b = 8'd117;  #10 
a = 8'd62; b = 8'd118;  #10 
a = 8'd62; b = 8'd119;  #10 
a = 8'd62; b = 8'd120;  #10 
a = 8'd62; b = 8'd121;  #10 
a = 8'd62; b = 8'd122;  #10 
a = 8'd62; b = 8'd123;  #10 
a = 8'd62; b = 8'd124;  #10 
a = 8'd62; b = 8'd125;  #10 
a = 8'd62; b = 8'd126;  #10 
a = 8'd62; b = 8'd127;  #10 
a = 8'd62; b = 8'd128;  #10 
a = 8'd62; b = 8'd129;  #10 
a = 8'd62; b = 8'd130;  #10 
a = 8'd62; b = 8'd131;  #10 
a = 8'd62; b = 8'd132;  #10 
a = 8'd62; b = 8'd133;  #10 
a = 8'd62; b = 8'd134;  #10 
a = 8'd62; b = 8'd135;  #10 
a = 8'd62; b = 8'd136;  #10 
a = 8'd62; b = 8'd137;  #10 
a = 8'd62; b = 8'd138;  #10 
a = 8'd62; b = 8'd139;  #10 
a = 8'd62; b = 8'd140;  #10 
a = 8'd62; b = 8'd141;  #10 
a = 8'd62; b = 8'd142;  #10 
a = 8'd62; b = 8'd143;  #10 
a = 8'd62; b = 8'd144;  #10 
a = 8'd62; b = 8'd145;  #10 
a = 8'd62; b = 8'd146;  #10 
a = 8'd62; b = 8'd147;  #10 
a = 8'd62; b = 8'd148;  #10 
a = 8'd62; b = 8'd149;  #10 
a = 8'd62; b = 8'd150;  #10 
a = 8'd62; b = 8'd151;  #10 
a = 8'd62; b = 8'd152;  #10 
a = 8'd62; b = 8'd153;  #10 
a = 8'd62; b = 8'd154;  #10 
a = 8'd62; b = 8'd155;  #10 
a = 8'd62; b = 8'd156;  #10 
a = 8'd62; b = 8'd157;  #10 
a = 8'd62; b = 8'd158;  #10 
a = 8'd62; b = 8'd159;  #10 
a = 8'd62; b = 8'd160;  #10 
a = 8'd62; b = 8'd161;  #10 
a = 8'd62; b = 8'd162;  #10 
a = 8'd62; b = 8'd163;  #10 
a = 8'd62; b = 8'd164;  #10 
a = 8'd62; b = 8'd165;  #10 
a = 8'd62; b = 8'd166;  #10 
a = 8'd62; b = 8'd167;  #10 
a = 8'd62; b = 8'd168;  #10 
a = 8'd62; b = 8'd169;  #10 
a = 8'd62; b = 8'd170;  #10 
a = 8'd62; b = 8'd171;  #10 
a = 8'd62; b = 8'd172;  #10 
a = 8'd62; b = 8'd173;  #10 
a = 8'd62; b = 8'd174;  #10 
a = 8'd62; b = 8'd175;  #10 
a = 8'd62; b = 8'd176;  #10 
a = 8'd62; b = 8'd177;  #10 
a = 8'd62; b = 8'd178;  #10 
a = 8'd62; b = 8'd179;  #10 
a = 8'd62; b = 8'd180;  #10 
a = 8'd62; b = 8'd181;  #10 
a = 8'd62; b = 8'd182;  #10 
a = 8'd62; b = 8'd183;  #10 
a = 8'd62; b = 8'd184;  #10 
a = 8'd62; b = 8'd185;  #10 
a = 8'd62; b = 8'd186;  #10 
a = 8'd62; b = 8'd187;  #10 
a = 8'd62; b = 8'd188;  #10 
a = 8'd62; b = 8'd189;  #10 
a = 8'd62; b = 8'd190;  #10 
a = 8'd62; b = 8'd191;  #10 
a = 8'd62; b = 8'd192;  #10 
a = 8'd62; b = 8'd193;  #10 
a = 8'd62; b = 8'd194;  #10 
a = 8'd62; b = 8'd195;  #10 
a = 8'd62; b = 8'd196;  #10 
a = 8'd62; b = 8'd197;  #10 
a = 8'd62; b = 8'd198;  #10 
a = 8'd62; b = 8'd199;  #10 
a = 8'd62; b = 8'd200;  #10 
a = 8'd62; b = 8'd201;  #10 
a = 8'd62; b = 8'd202;  #10 
a = 8'd62; b = 8'd203;  #10 
a = 8'd62; b = 8'd204;  #10 
a = 8'd62; b = 8'd205;  #10 
a = 8'd62; b = 8'd206;  #10 
a = 8'd62; b = 8'd207;  #10 
a = 8'd62; b = 8'd208;  #10 
a = 8'd62; b = 8'd209;  #10 
a = 8'd62; b = 8'd210;  #10 
a = 8'd62; b = 8'd211;  #10 
a = 8'd62; b = 8'd212;  #10 
a = 8'd62; b = 8'd213;  #10 
a = 8'd62; b = 8'd214;  #10 
a = 8'd62; b = 8'd215;  #10 
a = 8'd62; b = 8'd216;  #10 
a = 8'd62; b = 8'd217;  #10 
a = 8'd62; b = 8'd218;  #10 
a = 8'd62; b = 8'd219;  #10 
a = 8'd62; b = 8'd220;  #10 
a = 8'd62; b = 8'd221;  #10 
a = 8'd62; b = 8'd222;  #10 
a = 8'd62; b = 8'd223;  #10 
a = 8'd62; b = 8'd224;  #10 
a = 8'd62; b = 8'd225;  #10 
a = 8'd62; b = 8'd226;  #10 
a = 8'd62; b = 8'd227;  #10 
a = 8'd62; b = 8'd228;  #10 
a = 8'd62; b = 8'd229;  #10 
a = 8'd62; b = 8'd230;  #10 
a = 8'd62; b = 8'd231;  #10 
a = 8'd62; b = 8'd232;  #10 
a = 8'd62; b = 8'd233;  #10 
a = 8'd62; b = 8'd234;  #10 
a = 8'd62; b = 8'd235;  #10 
a = 8'd62; b = 8'd236;  #10 
a = 8'd62; b = 8'd237;  #10 
a = 8'd62; b = 8'd238;  #10 
a = 8'd62; b = 8'd239;  #10 
a = 8'd62; b = 8'd240;  #10 
a = 8'd62; b = 8'd241;  #10 
a = 8'd62; b = 8'd242;  #10 
a = 8'd62; b = 8'd243;  #10 
a = 8'd62; b = 8'd244;  #10 
a = 8'd62; b = 8'd245;  #10 
a = 8'd62; b = 8'd246;  #10 
a = 8'd62; b = 8'd247;  #10 
a = 8'd62; b = 8'd248;  #10 
a = 8'd62; b = 8'd249;  #10 
a = 8'd62; b = 8'd250;  #10 
a = 8'd62; b = 8'd251;  #10 
a = 8'd62; b = 8'd252;  #10 
a = 8'd62; b = 8'd253;  #10 
a = 8'd62; b = 8'd254;  #10 
a = 8'd62; b = 8'd255;  #10 
a = 8'd63; b = 8'd0;  #10 
a = 8'd63; b = 8'd1;  #10 
a = 8'd63; b = 8'd2;  #10 
a = 8'd63; b = 8'd3;  #10 
a = 8'd63; b = 8'd4;  #10 
a = 8'd63; b = 8'd5;  #10 
a = 8'd63; b = 8'd6;  #10 
a = 8'd63; b = 8'd7;  #10 
a = 8'd63; b = 8'd8;  #10 
a = 8'd63; b = 8'd9;  #10 
a = 8'd63; b = 8'd10;  #10 
a = 8'd63; b = 8'd11;  #10 
a = 8'd63; b = 8'd12;  #10 
a = 8'd63; b = 8'd13;  #10 
a = 8'd63; b = 8'd14;  #10 
a = 8'd63; b = 8'd15;  #10 
a = 8'd63; b = 8'd16;  #10 
a = 8'd63; b = 8'd17;  #10 
a = 8'd63; b = 8'd18;  #10 
a = 8'd63; b = 8'd19;  #10 
a = 8'd63; b = 8'd20;  #10 
a = 8'd63; b = 8'd21;  #10 
a = 8'd63; b = 8'd22;  #10 
a = 8'd63; b = 8'd23;  #10 
a = 8'd63; b = 8'd24;  #10 
a = 8'd63; b = 8'd25;  #10 
a = 8'd63; b = 8'd26;  #10 
a = 8'd63; b = 8'd27;  #10 
a = 8'd63; b = 8'd28;  #10 
a = 8'd63; b = 8'd29;  #10 
a = 8'd63; b = 8'd30;  #10 
a = 8'd63; b = 8'd31;  #10 
a = 8'd63; b = 8'd32;  #10 
a = 8'd63; b = 8'd33;  #10 
a = 8'd63; b = 8'd34;  #10 
a = 8'd63; b = 8'd35;  #10 
a = 8'd63; b = 8'd36;  #10 
a = 8'd63; b = 8'd37;  #10 
a = 8'd63; b = 8'd38;  #10 
a = 8'd63; b = 8'd39;  #10 
a = 8'd63; b = 8'd40;  #10 
a = 8'd63; b = 8'd41;  #10 
a = 8'd63; b = 8'd42;  #10 
a = 8'd63; b = 8'd43;  #10 
a = 8'd63; b = 8'd44;  #10 
a = 8'd63; b = 8'd45;  #10 
a = 8'd63; b = 8'd46;  #10 
a = 8'd63; b = 8'd47;  #10 
a = 8'd63; b = 8'd48;  #10 
a = 8'd63; b = 8'd49;  #10 
a = 8'd63; b = 8'd50;  #10 
a = 8'd63; b = 8'd51;  #10 
a = 8'd63; b = 8'd52;  #10 
a = 8'd63; b = 8'd53;  #10 
a = 8'd63; b = 8'd54;  #10 
a = 8'd63; b = 8'd55;  #10 
a = 8'd63; b = 8'd56;  #10 
a = 8'd63; b = 8'd57;  #10 
a = 8'd63; b = 8'd58;  #10 
a = 8'd63; b = 8'd59;  #10 
a = 8'd63; b = 8'd60;  #10 
a = 8'd63; b = 8'd61;  #10 
a = 8'd63; b = 8'd62;  #10 
a = 8'd63; b = 8'd63;  #10 
a = 8'd63; b = 8'd64;  #10 
a = 8'd63; b = 8'd65;  #10 
a = 8'd63; b = 8'd66;  #10 
a = 8'd63; b = 8'd67;  #10 
a = 8'd63; b = 8'd68;  #10 
a = 8'd63; b = 8'd69;  #10 
a = 8'd63; b = 8'd70;  #10 
a = 8'd63; b = 8'd71;  #10 
a = 8'd63; b = 8'd72;  #10 
a = 8'd63; b = 8'd73;  #10 
a = 8'd63; b = 8'd74;  #10 
a = 8'd63; b = 8'd75;  #10 
a = 8'd63; b = 8'd76;  #10 
a = 8'd63; b = 8'd77;  #10 
a = 8'd63; b = 8'd78;  #10 
a = 8'd63; b = 8'd79;  #10 
a = 8'd63; b = 8'd80;  #10 
a = 8'd63; b = 8'd81;  #10 
a = 8'd63; b = 8'd82;  #10 
a = 8'd63; b = 8'd83;  #10 
a = 8'd63; b = 8'd84;  #10 
a = 8'd63; b = 8'd85;  #10 
a = 8'd63; b = 8'd86;  #10 
a = 8'd63; b = 8'd87;  #10 
a = 8'd63; b = 8'd88;  #10 
a = 8'd63; b = 8'd89;  #10 
a = 8'd63; b = 8'd90;  #10 
a = 8'd63; b = 8'd91;  #10 
a = 8'd63; b = 8'd92;  #10 
a = 8'd63; b = 8'd93;  #10 
a = 8'd63; b = 8'd94;  #10 
a = 8'd63; b = 8'd95;  #10 
a = 8'd63; b = 8'd96;  #10 
a = 8'd63; b = 8'd97;  #10 
a = 8'd63; b = 8'd98;  #10 
a = 8'd63; b = 8'd99;  #10 
a = 8'd63; b = 8'd100;  #10 
a = 8'd63; b = 8'd101;  #10 
a = 8'd63; b = 8'd102;  #10 
a = 8'd63; b = 8'd103;  #10 
a = 8'd63; b = 8'd104;  #10 
a = 8'd63; b = 8'd105;  #10 
a = 8'd63; b = 8'd106;  #10 
a = 8'd63; b = 8'd107;  #10 
a = 8'd63; b = 8'd108;  #10 
a = 8'd63; b = 8'd109;  #10 
a = 8'd63; b = 8'd110;  #10 
a = 8'd63; b = 8'd111;  #10 
a = 8'd63; b = 8'd112;  #10 
a = 8'd63; b = 8'd113;  #10 
a = 8'd63; b = 8'd114;  #10 
a = 8'd63; b = 8'd115;  #10 
a = 8'd63; b = 8'd116;  #10 
a = 8'd63; b = 8'd117;  #10 
a = 8'd63; b = 8'd118;  #10 
a = 8'd63; b = 8'd119;  #10 
a = 8'd63; b = 8'd120;  #10 
a = 8'd63; b = 8'd121;  #10 
a = 8'd63; b = 8'd122;  #10 
a = 8'd63; b = 8'd123;  #10 
a = 8'd63; b = 8'd124;  #10 
a = 8'd63; b = 8'd125;  #10 
a = 8'd63; b = 8'd126;  #10 
a = 8'd63; b = 8'd127;  #10 
a = 8'd63; b = 8'd128;  #10 
a = 8'd63; b = 8'd129;  #10 
a = 8'd63; b = 8'd130;  #10 
a = 8'd63; b = 8'd131;  #10 
a = 8'd63; b = 8'd132;  #10 
a = 8'd63; b = 8'd133;  #10 
a = 8'd63; b = 8'd134;  #10 
a = 8'd63; b = 8'd135;  #10 
a = 8'd63; b = 8'd136;  #10 
a = 8'd63; b = 8'd137;  #10 
a = 8'd63; b = 8'd138;  #10 
a = 8'd63; b = 8'd139;  #10 
a = 8'd63; b = 8'd140;  #10 
a = 8'd63; b = 8'd141;  #10 
a = 8'd63; b = 8'd142;  #10 
a = 8'd63; b = 8'd143;  #10 
a = 8'd63; b = 8'd144;  #10 
a = 8'd63; b = 8'd145;  #10 
a = 8'd63; b = 8'd146;  #10 
a = 8'd63; b = 8'd147;  #10 
a = 8'd63; b = 8'd148;  #10 
a = 8'd63; b = 8'd149;  #10 
a = 8'd63; b = 8'd150;  #10 
a = 8'd63; b = 8'd151;  #10 
a = 8'd63; b = 8'd152;  #10 
a = 8'd63; b = 8'd153;  #10 
a = 8'd63; b = 8'd154;  #10 
a = 8'd63; b = 8'd155;  #10 
a = 8'd63; b = 8'd156;  #10 
a = 8'd63; b = 8'd157;  #10 
a = 8'd63; b = 8'd158;  #10 
a = 8'd63; b = 8'd159;  #10 
a = 8'd63; b = 8'd160;  #10 
a = 8'd63; b = 8'd161;  #10 
a = 8'd63; b = 8'd162;  #10 
a = 8'd63; b = 8'd163;  #10 
a = 8'd63; b = 8'd164;  #10 
a = 8'd63; b = 8'd165;  #10 
a = 8'd63; b = 8'd166;  #10 
a = 8'd63; b = 8'd167;  #10 
a = 8'd63; b = 8'd168;  #10 
a = 8'd63; b = 8'd169;  #10 
a = 8'd63; b = 8'd170;  #10 
a = 8'd63; b = 8'd171;  #10 
a = 8'd63; b = 8'd172;  #10 
a = 8'd63; b = 8'd173;  #10 
a = 8'd63; b = 8'd174;  #10 
a = 8'd63; b = 8'd175;  #10 
a = 8'd63; b = 8'd176;  #10 
a = 8'd63; b = 8'd177;  #10 
a = 8'd63; b = 8'd178;  #10 
a = 8'd63; b = 8'd179;  #10 
a = 8'd63; b = 8'd180;  #10 
a = 8'd63; b = 8'd181;  #10 
a = 8'd63; b = 8'd182;  #10 
a = 8'd63; b = 8'd183;  #10 
a = 8'd63; b = 8'd184;  #10 
a = 8'd63; b = 8'd185;  #10 
a = 8'd63; b = 8'd186;  #10 
a = 8'd63; b = 8'd187;  #10 
a = 8'd63; b = 8'd188;  #10 
a = 8'd63; b = 8'd189;  #10 
a = 8'd63; b = 8'd190;  #10 
a = 8'd63; b = 8'd191;  #10 
a = 8'd63; b = 8'd192;  #10 
a = 8'd63; b = 8'd193;  #10 
a = 8'd63; b = 8'd194;  #10 
a = 8'd63; b = 8'd195;  #10 
a = 8'd63; b = 8'd196;  #10 
a = 8'd63; b = 8'd197;  #10 
a = 8'd63; b = 8'd198;  #10 
a = 8'd63; b = 8'd199;  #10 
a = 8'd63; b = 8'd200;  #10 
a = 8'd63; b = 8'd201;  #10 
a = 8'd63; b = 8'd202;  #10 
a = 8'd63; b = 8'd203;  #10 
a = 8'd63; b = 8'd204;  #10 
a = 8'd63; b = 8'd205;  #10 
a = 8'd63; b = 8'd206;  #10 
a = 8'd63; b = 8'd207;  #10 
a = 8'd63; b = 8'd208;  #10 
a = 8'd63; b = 8'd209;  #10 
a = 8'd63; b = 8'd210;  #10 
a = 8'd63; b = 8'd211;  #10 
a = 8'd63; b = 8'd212;  #10 
a = 8'd63; b = 8'd213;  #10 
a = 8'd63; b = 8'd214;  #10 
a = 8'd63; b = 8'd215;  #10 
a = 8'd63; b = 8'd216;  #10 
a = 8'd63; b = 8'd217;  #10 
a = 8'd63; b = 8'd218;  #10 
a = 8'd63; b = 8'd219;  #10 
a = 8'd63; b = 8'd220;  #10 
a = 8'd63; b = 8'd221;  #10 
a = 8'd63; b = 8'd222;  #10 
a = 8'd63; b = 8'd223;  #10 
a = 8'd63; b = 8'd224;  #10 
a = 8'd63; b = 8'd225;  #10 
a = 8'd63; b = 8'd226;  #10 
a = 8'd63; b = 8'd227;  #10 
a = 8'd63; b = 8'd228;  #10 
a = 8'd63; b = 8'd229;  #10 
a = 8'd63; b = 8'd230;  #10 
a = 8'd63; b = 8'd231;  #10 
a = 8'd63; b = 8'd232;  #10 
a = 8'd63; b = 8'd233;  #10 
a = 8'd63; b = 8'd234;  #10 
a = 8'd63; b = 8'd235;  #10 
a = 8'd63; b = 8'd236;  #10 
a = 8'd63; b = 8'd237;  #10 
a = 8'd63; b = 8'd238;  #10 
a = 8'd63; b = 8'd239;  #10 
a = 8'd63; b = 8'd240;  #10 
a = 8'd63; b = 8'd241;  #10 
a = 8'd63; b = 8'd242;  #10 
a = 8'd63; b = 8'd243;  #10 
a = 8'd63; b = 8'd244;  #10 
a = 8'd63; b = 8'd245;  #10 
a = 8'd63; b = 8'd246;  #10 
a = 8'd63; b = 8'd247;  #10 
a = 8'd63; b = 8'd248;  #10 
a = 8'd63; b = 8'd249;  #10 
a = 8'd63; b = 8'd250;  #10 
a = 8'd63; b = 8'd251;  #10 
a = 8'd63; b = 8'd252;  #10 
a = 8'd63; b = 8'd253;  #10 
a = 8'd63; b = 8'd254;  #10 
a = 8'd63; b = 8'd255;  #10 
a = 8'd64; b = 8'd0;  #10 
a = 8'd64; b = 8'd1;  #10 
a = 8'd64; b = 8'd2;  #10 
a = 8'd64; b = 8'd3;  #10 
a = 8'd64; b = 8'd4;  #10 
a = 8'd64; b = 8'd5;  #10 
a = 8'd64; b = 8'd6;  #10 
a = 8'd64; b = 8'd7;  #10 
a = 8'd64; b = 8'd8;  #10 
a = 8'd64; b = 8'd9;  #10 
a = 8'd64; b = 8'd10;  #10 
a = 8'd64; b = 8'd11;  #10 
a = 8'd64; b = 8'd12;  #10 
a = 8'd64; b = 8'd13;  #10 
a = 8'd64; b = 8'd14;  #10 
a = 8'd64; b = 8'd15;  #10 
a = 8'd64; b = 8'd16;  #10 
a = 8'd64; b = 8'd17;  #10 
a = 8'd64; b = 8'd18;  #10 
a = 8'd64; b = 8'd19;  #10 
a = 8'd64; b = 8'd20;  #10 
a = 8'd64; b = 8'd21;  #10 
a = 8'd64; b = 8'd22;  #10 
a = 8'd64; b = 8'd23;  #10 
a = 8'd64; b = 8'd24;  #10 
a = 8'd64; b = 8'd25;  #10 
a = 8'd64; b = 8'd26;  #10 
a = 8'd64; b = 8'd27;  #10 
a = 8'd64; b = 8'd28;  #10 
a = 8'd64; b = 8'd29;  #10 
a = 8'd64; b = 8'd30;  #10 
a = 8'd64; b = 8'd31;  #10 
a = 8'd64; b = 8'd32;  #10 
a = 8'd64; b = 8'd33;  #10 
a = 8'd64; b = 8'd34;  #10 
a = 8'd64; b = 8'd35;  #10 
a = 8'd64; b = 8'd36;  #10 
a = 8'd64; b = 8'd37;  #10 
a = 8'd64; b = 8'd38;  #10 
a = 8'd64; b = 8'd39;  #10 
a = 8'd64; b = 8'd40;  #10 
a = 8'd64; b = 8'd41;  #10 
a = 8'd64; b = 8'd42;  #10 
a = 8'd64; b = 8'd43;  #10 
a = 8'd64; b = 8'd44;  #10 
a = 8'd64; b = 8'd45;  #10 
a = 8'd64; b = 8'd46;  #10 
a = 8'd64; b = 8'd47;  #10 
a = 8'd64; b = 8'd48;  #10 
a = 8'd64; b = 8'd49;  #10 
a = 8'd64; b = 8'd50;  #10 
a = 8'd64; b = 8'd51;  #10 
a = 8'd64; b = 8'd52;  #10 
a = 8'd64; b = 8'd53;  #10 
a = 8'd64; b = 8'd54;  #10 
a = 8'd64; b = 8'd55;  #10 
a = 8'd64; b = 8'd56;  #10 
a = 8'd64; b = 8'd57;  #10 
a = 8'd64; b = 8'd58;  #10 
a = 8'd64; b = 8'd59;  #10 
a = 8'd64; b = 8'd60;  #10 
a = 8'd64; b = 8'd61;  #10 
a = 8'd64; b = 8'd62;  #10 
a = 8'd64; b = 8'd63;  #10 
a = 8'd64; b = 8'd64;  #10 
a = 8'd64; b = 8'd65;  #10 
a = 8'd64; b = 8'd66;  #10 
a = 8'd64; b = 8'd67;  #10 
a = 8'd64; b = 8'd68;  #10 
a = 8'd64; b = 8'd69;  #10 
a = 8'd64; b = 8'd70;  #10 
a = 8'd64; b = 8'd71;  #10 
a = 8'd64; b = 8'd72;  #10 
a = 8'd64; b = 8'd73;  #10 
a = 8'd64; b = 8'd74;  #10 
a = 8'd64; b = 8'd75;  #10 
a = 8'd64; b = 8'd76;  #10 
a = 8'd64; b = 8'd77;  #10 
a = 8'd64; b = 8'd78;  #10 
a = 8'd64; b = 8'd79;  #10 
a = 8'd64; b = 8'd80;  #10 
a = 8'd64; b = 8'd81;  #10 
a = 8'd64; b = 8'd82;  #10 
a = 8'd64; b = 8'd83;  #10 
a = 8'd64; b = 8'd84;  #10 
a = 8'd64; b = 8'd85;  #10 
a = 8'd64; b = 8'd86;  #10 
a = 8'd64; b = 8'd87;  #10 
a = 8'd64; b = 8'd88;  #10 
a = 8'd64; b = 8'd89;  #10 
a = 8'd64; b = 8'd90;  #10 
a = 8'd64; b = 8'd91;  #10 
a = 8'd64; b = 8'd92;  #10 
a = 8'd64; b = 8'd93;  #10 
a = 8'd64; b = 8'd94;  #10 
a = 8'd64; b = 8'd95;  #10 
a = 8'd64; b = 8'd96;  #10 
a = 8'd64; b = 8'd97;  #10 
a = 8'd64; b = 8'd98;  #10 
a = 8'd64; b = 8'd99;  #10 
a = 8'd64; b = 8'd100;  #10 
a = 8'd64; b = 8'd101;  #10 
a = 8'd64; b = 8'd102;  #10 
a = 8'd64; b = 8'd103;  #10 
a = 8'd64; b = 8'd104;  #10 
a = 8'd64; b = 8'd105;  #10 
a = 8'd64; b = 8'd106;  #10 
a = 8'd64; b = 8'd107;  #10 
a = 8'd64; b = 8'd108;  #10 
a = 8'd64; b = 8'd109;  #10 
a = 8'd64; b = 8'd110;  #10 
a = 8'd64; b = 8'd111;  #10 
a = 8'd64; b = 8'd112;  #10 
a = 8'd64; b = 8'd113;  #10 
a = 8'd64; b = 8'd114;  #10 
a = 8'd64; b = 8'd115;  #10 
a = 8'd64; b = 8'd116;  #10 
a = 8'd64; b = 8'd117;  #10 
a = 8'd64; b = 8'd118;  #10 
a = 8'd64; b = 8'd119;  #10 
a = 8'd64; b = 8'd120;  #10 
a = 8'd64; b = 8'd121;  #10 
a = 8'd64; b = 8'd122;  #10 
a = 8'd64; b = 8'd123;  #10 
a = 8'd64; b = 8'd124;  #10 
a = 8'd64; b = 8'd125;  #10 
a = 8'd64; b = 8'd126;  #10 
a = 8'd64; b = 8'd127;  #10 
a = 8'd64; b = 8'd128;  #10 
a = 8'd64; b = 8'd129;  #10 
a = 8'd64; b = 8'd130;  #10 
a = 8'd64; b = 8'd131;  #10 
a = 8'd64; b = 8'd132;  #10 
a = 8'd64; b = 8'd133;  #10 
a = 8'd64; b = 8'd134;  #10 
a = 8'd64; b = 8'd135;  #10 
a = 8'd64; b = 8'd136;  #10 
a = 8'd64; b = 8'd137;  #10 
a = 8'd64; b = 8'd138;  #10 
a = 8'd64; b = 8'd139;  #10 
a = 8'd64; b = 8'd140;  #10 
a = 8'd64; b = 8'd141;  #10 
a = 8'd64; b = 8'd142;  #10 
a = 8'd64; b = 8'd143;  #10 
a = 8'd64; b = 8'd144;  #10 
a = 8'd64; b = 8'd145;  #10 
a = 8'd64; b = 8'd146;  #10 
a = 8'd64; b = 8'd147;  #10 
a = 8'd64; b = 8'd148;  #10 
a = 8'd64; b = 8'd149;  #10 
a = 8'd64; b = 8'd150;  #10 
a = 8'd64; b = 8'd151;  #10 
a = 8'd64; b = 8'd152;  #10 
a = 8'd64; b = 8'd153;  #10 
a = 8'd64; b = 8'd154;  #10 
a = 8'd64; b = 8'd155;  #10 
a = 8'd64; b = 8'd156;  #10 
a = 8'd64; b = 8'd157;  #10 
a = 8'd64; b = 8'd158;  #10 
a = 8'd64; b = 8'd159;  #10 
a = 8'd64; b = 8'd160;  #10 
a = 8'd64; b = 8'd161;  #10 
a = 8'd64; b = 8'd162;  #10 
a = 8'd64; b = 8'd163;  #10 
a = 8'd64; b = 8'd164;  #10 
a = 8'd64; b = 8'd165;  #10 
a = 8'd64; b = 8'd166;  #10 
a = 8'd64; b = 8'd167;  #10 
a = 8'd64; b = 8'd168;  #10 
a = 8'd64; b = 8'd169;  #10 
a = 8'd64; b = 8'd170;  #10 
a = 8'd64; b = 8'd171;  #10 
a = 8'd64; b = 8'd172;  #10 
a = 8'd64; b = 8'd173;  #10 
a = 8'd64; b = 8'd174;  #10 
a = 8'd64; b = 8'd175;  #10 
a = 8'd64; b = 8'd176;  #10 
a = 8'd64; b = 8'd177;  #10 
a = 8'd64; b = 8'd178;  #10 
a = 8'd64; b = 8'd179;  #10 
a = 8'd64; b = 8'd180;  #10 
a = 8'd64; b = 8'd181;  #10 
a = 8'd64; b = 8'd182;  #10 
a = 8'd64; b = 8'd183;  #10 
a = 8'd64; b = 8'd184;  #10 
a = 8'd64; b = 8'd185;  #10 
a = 8'd64; b = 8'd186;  #10 
a = 8'd64; b = 8'd187;  #10 
a = 8'd64; b = 8'd188;  #10 
a = 8'd64; b = 8'd189;  #10 
a = 8'd64; b = 8'd190;  #10 
a = 8'd64; b = 8'd191;  #10 
a = 8'd64; b = 8'd192;  #10 
a = 8'd64; b = 8'd193;  #10 
a = 8'd64; b = 8'd194;  #10 
a = 8'd64; b = 8'd195;  #10 
a = 8'd64; b = 8'd196;  #10 
a = 8'd64; b = 8'd197;  #10 
a = 8'd64; b = 8'd198;  #10 
a = 8'd64; b = 8'd199;  #10 
a = 8'd64; b = 8'd200;  #10 
a = 8'd64; b = 8'd201;  #10 
a = 8'd64; b = 8'd202;  #10 
a = 8'd64; b = 8'd203;  #10 
a = 8'd64; b = 8'd204;  #10 
a = 8'd64; b = 8'd205;  #10 
a = 8'd64; b = 8'd206;  #10 
a = 8'd64; b = 8'd207;  #10 
a = 8'd64; b = 8'd208;  #10 
a = 8'd64; b = 8'd209;  #10 
a = 8'd64; b = 8'd210;  #10 
a = 8'd64; b = 8'd211;  #10 
a = 8'd64; b = 8'd212;  #10 
a = 8'd64; b = 8'd213;  #10 
a = 8'd64; b = 8'd214;  #10 
a = 8'd64; b = 8'd215;  #10 
a = 8'd64; b = 8'd216;  #10 
a = 8'd64; b = 8'd217;  #10 
a = 8'd64; b = 8'd218;  #10 
a = 8'd64; b = 8'd219;  #10 
a = 8'd64; b = 8'd220;  #10 
a = 8'd64; b = 8'd221;  #10 
a = 8'd64; b = 8'd222;  #10 
a = 8'd64; b = 8'd223;  #10 
a = 8'd64; b = 8'd224;  #10 
a = 8'd64; b = 8'd225;  #10 
a = 8'd64; b = 8'd226;  #10 
a = 8'd64; b = 8'd227;  #10 
a = 8'd64; b = 8'd228;  #10 
a = 8'd64; b = 8'd229;  #10 
a = 8'd64; b = 8'd230;  #10 
a = 8'd64; b = 8'd231;  #10 
a = 8'd64; b = 8'd232;  #10 
a = 8'd64; b = 8'd233;  #10 
a = 8'd64; b = 8'd234;  #10 
a = 8'd64; b = 8'd235;  #10 
a = 8'd64; b = 8'd236;  #10 
a = 8'd64; b = 8'd237;  #10 
a = 8'd64; b = 8'd238;  #10 
a = 8'd64; b = 8'd239;  #10 
a = 8'd64; b = 8'd240;  #10 
a = 8'd64; b = 8'd241;  #10 
a = 8'd64; b = 8'd242;  #10 
a = 8'd64; b = 8'd243;  #10 
a = 8'd64; b = 8'd244;  #10 
a = 8'd64; b = 8'd245;  #10 
a = 8'd64; b = 8'd246;  #10 
a = 8'd64; b = 8'd247;  #10 
a = 8'd64; b = 8'd248;  #10 
a = 8'd64; b = 8'd249;  #10 
a = 8'd64; b = 8'd250;  #10 
a = 8'd64; b = 8'd251;  #10 
a = 8'd64; b = 8'd252;  #10 
a = 8'd64; b = 8'd253;  #10 
a = 8'd64; b = 8'd254;  #10 
a = 8'd64; b = 8'd255;  #10 
a = 8'd65; b = 8'd0;  #10 
a = 8'd65; b = 8'd1;  #10 
a = 8'd65; b = 8'd2;  #10 
a = 8'd65; b = 8'd3;  #10 
a = 8'd65; b = 8'd4;  #10 
a = 8'd65; b = 8'd5;  #10 
a = 8'd65; b = 8'd6;  #10 
a = 8'd65; b = 8'd7;  #10 
a = 8'd65; b = 8'd8;  #10 
a = 8'd65; b = 8'd9;  #10 
a = 8'd65; b = 8'd10;  #10 
a = 8'd65; b = 8'd11;  #10 
a = 8'd65; b = 8'd12;  #10 
a = 8'd65; b = 8'd13;  #10 
a = 8'd65; b = 8'd14;  #10 
a = 8'd65; b = 8'd15;  #10 
a = 8'd65; b = 8'd16;  #10 
a = 8'd65; b = 8'd17;  #10 
a = 8'd65; b = 8'd18;  #10 
a = 8'd65; b = 8'd19;  #10 
a = 8'd65; b = 8'd20;  #10 
a = 8'd65; b = 8'd21;  #10 
a = 8'd65; b = 8'd22;  #10 
a = 8'd65; b = 8'd23;  #10 
a = 8'd65; b = 8'd24;  #10 
a = 8'd65; b = 8'd25;  #10 
a = 8'd65; b = 8'd26;  #10 
a = 8'd65; b = 8'd27;  #10 
a = 8'd65; b = 8'd28;  #10 
a = 8'd65; b = 8'd29;  #10 
a = 8'd65; b = 8'd30;  #10 
a = 8'd65; b = 8'd31;  #10 
a = 8'd65; b = 8'd32;  #10 
a = 8'd65; b = 8'd33;  #10 
a = 8'd65; b = 8'd34;  #10 
a = 8'd65; b = 8'd35;  #10 
a = 8'd65; b = 8'd36;  #10 
a = 8'd65; b = 8'd37;  #10 
a = 8'd65; b = 8'd38;  #10 
a = 8'd65; b = 8'd39;  #10 
a = 8'd65; b = 8'd40;  #10 
a = 8'd65; b = 8'd41;  #10 
a = 8'd65; b = 8'd42;  #10 
a = 8'd65; b = 8'd43;  #10 
a = 8'd65; b = 8'd44;  #10 
a = 8'd65; b = 8'd45;  #10 
a = 8'd65; b = 8'd46;  #10 
a = 8'd65; b = 8'd47;  #10 
a = 8'd65; b = 8'd48;  #10 
a = 8'd65; b = 8'd49;  #10 
a = 8'd65; b = 8'd50;  #10 
a = 8'd65; b = 8'd51;  #10 
a = 8'd65; b = 8'd52;  #10 
a = 8'd65; b = 8'd53;  #10 
a = 8'd65; b = 8'd54;  #10 
a = 8'd65; b = 8'd55;  #10 
a = 8'd65; b = 8'd56;  #10 
a = 8'd65; b = 8'd57;  #10 
a = 8'd65; b = 8'd58;  #10 
a = 8'd65; b = 8'd59;  #10 
a = 8'd65; b = 8'd60;  #10 
a = 8'd65; b = 8'd61;  #10 
a = 8'd65; b = 8'd62;  #10 
a = 8'd65; b = 8'd63;  #10 
a = 8'd65; b = 8'd64;  #10 
a = 8'd65; b = 8'd65;  #10 
a = 8'd65; b = 8'd66;  #10 
a = 8'd65; b = 8'd67;  #10 
a = 8'd65; b = 8'd68;  #10 
a = 8'd65; b = 8'd69;  #10 
a = 8'd65; b = 8'd70;  #10 
a = 8'd65; b = 8'd71;  #10 
a = 8'd65; b = 8'd72;  #10 
a = 8'd65; b = 8'd73;  #10 
a = 8'd65; b = 8'd74;  #10 
a = 8'd65; b = 8'd75;  #10 
a = 8'd65; b = 8'd76;  #10 
a = 8'd65; b = 8'd77;  #10 
a = 8'd65; b = 8'd78;  #10 
a = 8'd65; b = 8'd79;  #10 
a = 8'd65; b = 8'd80;  #10 
a = 8'd65; b = 8'd81;  #10 
a = 8'd65; b = 8'd82;  #10 
a = 8'd65; b = 8'd83;  #10 
a = 8'd65; b = 8'd84;  #10 
a = 8'd65; b = 8'd85;  #10 
a = 8'd65; b = 8'd86;  #10 
a = 8'd65; b = 8'd87;  #10 
a = 8'd65; b = 8'd88;  #10 
a = 8'd65; b = 8'd89;  #10 
a = 8'd65; b = 8'd90;  #10 
a = 8'd65; b = 8'd91;  #10 
a = 8'd65; b = 8'd92;  #10 
a = 8'd65; b = 8'd93;  #10 
a = 8'd65; b = 8'd94;  #10 
a = 8'd65; b = 8'd95;  #10 
a = 8'd65; b = 8'd96;  #10 
a = 8'd65; b = 8'd97;  #10 
a = 8'd65; b = 8'd98;  #10 
a = 8'd65; b = 8'd99;  #10 
a = 8'd65; b = 8'd100;  #10 
a = 8'd65; b = 8'd101;  #10 
a = 8'd65; b = 8'd102;  #10 
a = 8'd65; b = 8'd103;  #10 
a = 8'd65; b = 8'd104;  #10 
a = 8'd65; b = 8'd105;  #10 
a = 8'd65; b = 8'd106;  #10 
a = 8'd65; b = 8'd107;  #10 
a = 8'd65; b = 8'd108;  #10 
a = 8'd65; b = 8'd109;  #10 
a = 8'd65; b = 8'd110;  #10 
a = 8'd65; b = 8'd111;  #10 
a = 8'd65; b = 8'd112;  #10 
a = 8'd65; b = 8'd113;  #10 
a = 8'd65; b = 8'd114;  #10 
a = 8'd65; b = 8'd115;  #10 
a = 8'd65; b = 8'd116;  #10 
a = 8'd65; b = 8'd117;  #10 
a = 8'd65; b = 8'd118;  #10 
a = 8'd65; b = 8'd119;  #10 
a = 8'd65; b = 8'd120;  #10 
a = 8'd65; b = 8'd121;  #10 
a = 8'd65; b = 8'd122;  #10 
a = 8'd65; b = 8'd123;  #10 
a = 8'd65; b = 8'd124;  #10 
a = 8'd65; b = 8'd125;  #10 
a = 8'd65; b = 8'd126;  #10 
a = 8'd65; b = 8'd127;  #10 
a = 8'd65; b = 8'd128;  #10 
a = 8'd65; b = 8'd129;  #10 
a = 8'd65; b = 8'd130;  #10 
a = 8'd65; b = 8'd131;  #10 
a = 8'd65; b = 8'd132;  #10 
a = 8'd65; b = 8'd133;  #10 
a = 8'd65; b = 8'd134;  #10 
a = 8'd65; b = 8'd135;  #10 
a = 8'd65; b = 8'd136;  #10 
a = 8'd65; b = 8'd137;  #10 
a = 8'd65; b = 8'd138;  #10 
a = 8'd65; b = 8'd139;  #10 
a = 8'd65; b = 8'd140;  #10 
a = 8'd65; b = 8'd141;  #10 
a = 8'd65; b = 8'd142;  #10 
a = 8'd65; b = 8'd143;  #10 
a = 8'd65; b = 8'd144;  #10 
a = 8'd65; b = 8'd145;  #10 
a = 8'd65; b = 8'd146;  #10 
a = 8'd65; b = 8'd147;  #10 
a = 8'd65; b = 8'd148;  #10 
a = 8'd65; b = 8'd149;  #10 
a = 8'd65; b = 8'd150;  #10 
a = 8'd65; b = 8'd151;  #10 
a = 8'd65; b = 8'd152;  #10 
a = 8'd65; b = 8'd153;  #10 
a = 8'd65; b = 8'd154;  #10 
a = 8'd65; b = 8'd155;  #10 
a = 8'd65; b = 8'd156;  #10 
a = 8'd65; b = 8'd157;  #10 
a = 8'd65; b = 8'd158;  #10 
a = 8'd65; b = 8'd159;  #10 
a = 8'd65; b = 8'd160;  #10 
a = 8'd65; b = 8'd161;  #10 
a = 8'd65; b = 8'd162;  #10 
a = 8'd65; b = 8'd163;  #10 
a = 8'd65; b = 8'd164;  #10 
a = 8'd65; b = 8'd165;  #10 
a = 8'd65; b = 8'd166;  #10 
a = 8'd65; b = 8'd167;  #10 
a = 8'd65; b = 8'd168;  #10 
a = 8'd65; b = 8'd169;  #10 
a = 8'd65; b = 8'd170;  #10 
a = 8'd65; b = 8'd171;  #10 
a = 8'd65; b = 8'd172;  #10 
a = 8'd65; b = 8'd173;  #10 
a = 8'd65; b = 8'd174;  #10 
a = 8'd65; b = 8'd175;  #10 
a = 8'd65; b = 8'd176;  #10 
a = 8'd65; b = 8'd177;  #10 
a = 8'd65; b = 8'd178;  #10 
a = 8'd65; b = 8'd179;  #10 
a = 8'd65; b = 8'd180;  #10 
a = 8'd65; b = 8'd181;  #10 
a = 8'd65; b = 8'd182;  #10 
a = 8'd65; b = 8'd183;  #10 
a = 8'd65; b = 8'd184;  #10 
a = 8'd65; b = 8'd185;  #10 
a = 8'd65; b = 8'd186;  #10 
a = 8'd65; b = 8'd187;  #10 
a = 8'd65; b = 8'd188;  #10 
a = 8'd65; b = 8'd189;  #10 
a = 8'd65; b = 8'd190;  #10 
a = 8'd65; b = 8'd191;  #10 
a = 8'd65; b = 8'd192;  #10 
a = 8'd65; b = 8'd193;  #10 
a = 8'd65; b = 8'd194;  #10 
a = 8'd65; b = 8'd195;  #10 
a = 8'd65; b = 8'd196;  #10 
a = 8'd65; b = 8'd197;  #10 
a = 8'd65; b = 8'd198;  #10 
a = 8'd65; b = 8'd199;  #10 
a = 8'd65; b = 8'd200;  #10 
a = 8'd65; b = 8'd201;  #10 
a = 8'd65; b = 8'd202;  #10 
a = 8'd65; b = 8'd203;  #10 
a = 8'd65; b = 8'd204;  #10 
a = 8'd65; b = 8'd205;  #10 
a = 8'd65; b = 8'd206;  #10 
a = 8'd65; b = 8'd207;  #10 
a = 8'd65; b = 8'd208;  #10 
a = 8'd65; b = 8'd209;  #10 
a = 8'd65; b = 8'd210;  #10 
a = 8'd65; b = 8'd211;  #10 
a = 8'd65; b = 8'd212;  #10 
a = 8'd65; b = 8'd213;  #10 
a = 8'd65; b = 8'd214;  #10 
a = 8'd65; b = 8'd215;  #10 
a = 8'd65; b = 8'd216;  #10 
a = 8'd65; b = 8'd217;  #10 
a = 8'd65; b = 8'd218;  #10 
a = 8'd65; b = 8'd219;  #10 
a = 8'd65; b = 8'd220;  #10 
a = 8'd65; b = 8'd221;  #10 
a = 8'd65; b = 8'd222;  #10 
a = 8'd65; b = 8'd223;  #10 
a = 8'd65; b = 8'd224;  #10 
a = 8'd65; b = 8'd225;  #10 
a = 8'd65; b = 8'd226;  #10 
a = 8'd65; b = 8'd227;  #10 
a = 8'd65; b = 8'd228;  #10 
a = 8'd65; b = 8'd229;  #10 
a = 8'd65; b = 8'd230;  #10 
a = 8'd65; b = 8'd231;  #10 
a = 8'd65; b = 8'd232;  #10 
a = 8'd65; b = 8'd233;  #10 
a = 8'd65; b = 8'd234;  #10 
a = 8'd65; b = 8'd235;  #10 
a = 8'd65; b = 8'd236;  #10 
a = 8'd65; b = 8'd237;  #10 
a = 8'd65; b = 8'd238;  #10 
a = 8'd65; b = 8'd239;  #10 
a = 8'd65; b = 8'd240;  #10 
a = 8'd65; b = 8'd241;  #10 
a = 8'd65; b = 8'd242;  #10 
a = 8'd65; b = 8'd243;  #10 
a = 8'd65; b = 8'd244;  #10 
a = 8'd65; b = 8'd245;  #10 
a = 8'd65; b = 8'd246;  #10 
a = 8'd65; b = 8'd247;  #10 
a = 8'd65; b = 8'd248;  #10 
a = 8'd65; b = 8'd249;  #10 
a = 8'd65; b = 8'd250;  #10 
a = 8'd65; b = 8'd251;  #10 
a = 8'd65; b = 8'd252;  #10 
a = 8'd65; b = 8'd253;  #10 
a = 8'd65; b = 8'd254;  #10 
a = 8'd65; b = 8'd255;  #10 
a = 8'd66; b = 8'd0;  #10 
a = 8'd66; b = 8'd1;  #10 
a = 8'd66; b = 8'd2;  #10 
a = 8'd66; b = 8'd3;  #10 
a = 8'd66; b = 8'd4;  #10 
a = 8'd66; b = 8'd5;  #10 
a = 8'd66; b = 8'd6;  #10 
a = 8'd66; b = 8'd7;  #10 
a = 8'd66; b = 8'd8;  #10 
a = 8'd66; b = 8'd9;  #10 
a = 8'd66; b = 8'd10;  #10 
a = 8'd66; b = 8'd11;  #10 
a = 8'd66; b = 8'd12;  #10 
a = 8'd66; b = 8'd13;  #10 
a = 8'd66; b = 8'd14;  #10 
a = 8'd66; b = 8'd15;  #10 
a = 8'd66; b = 8'd16;  #10 
a = 8'd66; b = 8'd17;  #10 
a = 8'd66; b = 8'd18;  #10 
a = 8'd66; b = 8'd19;  #10 
a = 8'd66; b = 8'd20;  #10 
a = 8'd66; b = 8'd21;  #10 
a = 8'd66; b = 8'd22;  #10 
a = 8'd66; b = 8'd23;  #10 
a = 8'd66; b = 8'd24;  #10 
a = 8'd66; b = 8'd25;  #10 
a = 8'd66; b = 8'd26;  #10 
a = 8'd66; b = 8'd27;  #10 
a = 8'd66; b = 8'd28;  #10 
a = 8'd66; b = 8'd29;  #10 
a = 8'd66; b = 8'd30;  #10 
a = 8'd66; b = 8'd31;  #10 
a = 8'd66; b = 8'd32;  #10 
a = 8'd66; b = 8'd33;  #10 
a = 8'd66; b = 8'd34;  #10 
a = 8'd66; b = 8'd35;  #10 
a = 8'd66; b = 8'd36;  #10 
a = 8'd66; b = 8'd37;  #10 
a = 8'd66; b = 8'd38;  #10 
a = 8'd66; b = 8'd39;  #10 
a = 8'd66; b = 8'd40;  #10 
a = 8'd66; b = 8'd41;  #10 
a = 8'd66; b = 8'd42;  #10 
a = 8'd66; b = 8'd43;  #10 
a = 8'd66; b = 8'd44;  #10 
a = 8'd66; b = 8'd45;  #10 
a = 8'd66; b = 8'd46;  #10 
a = 8'd66; b = 8'd47;  #10 
a = 8'd66; b = 8'd48;  #10 
a = 8'd66; b = 8'd49;  #10 
a = 8'd66; b = 8'd50;  #10 
a = 8'd66; b = 8'd51;  #10 
a = 8'd66; b = 8'd52;  #10 
a = 8'd66; b = 8'd53;  #10 
a = 8'd66; b = 8'd54;  #10 
a = 8'd66; b = 8'd55;  #10 
a = 8'd66; b = 8'd56;  #10 
a = 8'd66; b = 8'd57;  #10 
a = 8'd66; b = 8'd58;  #10 
a = 8'd66; b = 8'd59;  #10 
a = 8'd66; b = 8'd60;  #10 
a = 8'd66; b = 8'd61;  #10 
a = 8'd66; b = 8'd62;  #10 
a = 8'd66; b = 8'd63;  #10 
a = 8'd66; b = 8'd64;  #10 
a = 8'd66; b = 8'd65;  #10 
a = 8'd66; b = 8'd66;  #10 
a = 8'd66; b = 8'd67;  #10 
a = 8'd66; b = 8'd68;  #10 
a = 8'd66; b = 8'd69;  #10 
a = 8'd66; b = 8'd70;  #10 
a = 8'd66; b = 8'd71;  #10 
a = 8'd66; b = 8'd72;  #10 
a = 8'd66; b = 8'd73;  #10 
a = 8'd66; b = 8'd74;  #10 
a = 8'd66; b = 8'd75;  #10 
a = 8'd66; b = 8'd76;  #10 
a = 8'd66; b = 8'd77;  #10 
a = 8'd66; b = 8'd78;  #10 
a = 8'd66; b = 8'd79;  #10 
a = 8'd66; b = 8'd80;  #10 
a = 8'd66; b = 8'd81;  #10 
a = 8'd66; b = 8'd82;  #10 
a = 8'd66; b = 8'd83;  #10 
a = 8'd66; b = 8'd84;  #10 
a = 8'd66; b = 8'd85;  #10 
a = 8'd66; b = 8'd86;  #10 
a = 8'd66; b = 8'd87;  #10 
a = 8'd66; b = 8'd88;  #10 
a = 8'd66; b = 8'd89;  #10 
a = 8'd66; b = 8'd90;  #10 
a = 8'd66; b = 8'd91;  #10 
a = 8'd66; b = 8'd92;  #10 
a = 8'd66; b = 8'd93;  #10 
a = 8'd66; b = 8'd94;  #10 
a = 8'd66; b = 8'd95;  #10 
a = 8'd66; b = 8'd96;  #10 
a = 8'd66; b = 8'd97;  #10 
a = 8'd66; b = 8'd98;  #10 
a = 8'd66; b = 8'd99;  #10 
a = 8'd66; b = 8'd100;  #10 
a = 8'd66; b = 8'd101;  #10 
a = 8'd66; b = 8'd102;  #10 
a = 8'd66; b = 8'd103;  #10 
a = 8'd66; b = 8'd104;  #10 
a = 8'd66; b = 8'd105;  #10 
a = 8'd66; b = 8'd106;  #10 
a = 8'd66; b = 8'd107;  #10 
a = 8'd66; b = 8'd108;  #10 
a = 8'd66; b = 8'd109;  #10 
a = 8'd66; b = 8'd110;  #10 
a = 8'd66; b = 8'd111;  #10 
a = 8'd66; b = 8'd112;  #10 
a = 8'd66; b = 8'd113;  #10 
a = 8'd66; b = 8'd114;  #10 
a = 8'd66; b = 8'd115;  #10 
a = 8'd66; b = 8'd116;  #10 
a = 8'd66; b = 8'd117;  #10 
a = 8'd66; b = 8'd118;  #10 
a = 8'd66; b = 8'd119;  #10 
a = 8'd66; b = 8'd120;  #10 
a = 8'd66; b = 8'd121;  #10 
a = 8'd66; b = 8'd122;  #10 
a = 8'd66; b = 8'd123;  #10 
a = 8'd66; b = 8'd124;  #10 
a = 8'd66; b = 8'd125;  #10 
a = 8'd66; b = 8'd126;  #10 
a = 8'd66; b = 8'd127;  #10 
a = 8'd66; b = 8'd128;  #10 
a = 8'd66; b = 8'd129;  #10 
a = 8'd66; b = 8'd130;  #10 
a = 8'd66; b = 8'd131;  #10 
a = 8'd66; b = 8'd132;  #10 
a = 8'd66; b = 8'd133;  #10 
a = 8'd66; b = 8'd134;  #10 
a = 8'd66; b = 8'd135;  #10 
a = 8'd66; b = 8'd136;  #10 
a = 8'd66; b = 8'd137;  #10 
a = 8'd66; b = 8'd138;  #10 
a = 8'd66; b = 8'd139;  #10 
a = 8'd66; b = 8'd140;  #10 
a = 8'd66; b = 8'd141;  #10 
a = 8'd66; b = 8'd142;  #10 
a = 8'd66; b = 8'd143;  #10 
a = 8'd66; b = 8'd144;  #10 
a = 8'd66; b = 8'd145;  #10 
a = 8'd66; b = 8'd146;  #10 
a = 8'd66; b = 8'd147;  #10 
a = 8'd66; b = 8'd148;  #10 
a = 8'd66; b = 8'd149;  #10 
a = 8'd66; b = 8'd150;  #10 
a = 8'd66; b = 8'd151;  #10 
a = 8'd66; b = 8'd152;  #10 
a = 8'd66; b = 8'd153;  #10 
a = 8'd66; b = 8'd154;  #10 
a = 8'd66; b = 8'd155;  #10 
a = 8'd66; b = 8'd156;  #10 
a = 8'd66; b = 8'd157;  #10 
a = 8'd66; b = 8'd158;  #10 
a = 8'd66; b = 8'd159;  #10 
a = 8'd66; b = 8'd160;  #10 
a = 8'd66; b = 8'd161;  #10 
a = 8'd66; b = 8'd162;  #10 
a = 8'd66; b = 8'd163;  #10 
a = 8'd66; b = 8'd164;  #10 
a = 8'd66; b = 8'd165;  #10 
a = 8'd66; b = 8'd166;  #10 
a = 8'd66; b = 8'd167;  #10 
a = 8'd66; b = 8'd168;  #10 
a = 8'd66; b = 8'd169;  #10 
a = 8'd66; b = 8'd170;  #10 
a = 8'd66; b = 8'd171;  #10 
a = 8'd66; b = 8'd172;  #10 
a = 8'd66; b = 8'd173;  #10 
a = 8'd66; b = 8'd174;  #10 
a = 8'd66; b = 8'd175;  #10 
a = 8'd66; b = 8'd176;  #10 
a = 8'd66; b = 8'd177;  #10 
a = 8'd66; b = 8'd178;  #10 
a = 8'd66; b = 8'd179;  #10 
a = 8'd66; b = 8'd180;  #10 
a = 8'd66; b = 8'd181;  #10 
a = 8'd66; b = 8'd182;  #10 
a = 8'd66; b = 8'd183;  #10 
a = 8'd66; b = 8'd184;  #10 
a = 8'd66; b = 8'd185;  #10 
a = 8'd66; b = 8'd186;  #10 
a = 8'd66; b = 8'd187;  #10 
a = 8'd66; b = 8'd188;  #10 
a = 8'd66; b = 8'd189;  #10 
a = 8'd66; b = 8'd190;  #10 
a = 8'd66; b = 8'd191;  #10 
a = 8'd66; b = 8'd192;  #10 
a = 8'd66; b = 8'd193;  #10 
a = 8'd66; b = 8'd194;  #10 
a = 8'd66; b = 8'd195;  #10 
a = 8'd66; b = 8'd196;  #10 
a = 8'd66; b = 8'd197;  #10 
a = 8'd66; b = 8'd198;  #10 
a = 8'd66; b = 8'd199;  #10 
a = 8'd66; b = 8'd200;  #10 
a = 8'd66; b = 8'd201;  #10 
a = 8'd66; b = 8'd202;  #10 
a = 8'd66; b = 8'd203;  #10 
a = 8'd66; b = 8'd204;  #10 
a = 8'd66; b = 8'd205;  #10 
a = 8'd66; b = 8'd206;  #10 
a = 8'd66; b = 8'd207;  #10 
a = 8'd66; b = 8'd208;  #10 
a = 8'd66; b = 8'd209;  #10 
a = 8'd66; b = 8'd210;  #10 
a = 8'd66; b = 8'd211;  #10 
a = 8'd66; b = 8'd212;  #10 
a = 8'd66; b = 8'd213;  #10 
a = 8'd66; b = 8'd214;  #10 
a = 8'd66; b = 8'd215;  #10 
a = 8'd66; b = 8'd216;  #10 
a = 8'd66; b = 8'd217;  #10 
a = 8'd66; b = 8'd218;  #10 
a = 8'd66; b = 8'd219;  #10 
a = 8'd66; b = 8'd220;  #10 
a = 8'd66; b = 8'd221;  #10 
a = 8'd66; b = 8'd222;  #10 
a = 8'd66; b = 8'd223;  #10 
a = 8'd66; b = 8'd224;  #10 
a = 8'd66; b = 8'd225;  #10 
a = 8'd66; b = 8'd226;  #10 
a = 8'd66; b = 8'd227;  #10 
a = 8'd66; b = 8'd228;  #10 
a = 8'd66; b = 8'd229;  #10 
a = 8'd66; b = 8'd230;  #10 
a = 8'd66; b = 8'd231;  #10 
a = 8'd66; b = 8'd232;  #10 
a = 8'd66; b = 8'd233;  #10 
a = 8'd66; b = 8'd234;  #10 
a = 8'd66; b = 8'd235;  #10 
a = 8'd66; b = 8'd236;  #10 
a = 8'd66; b = 8'd237;  #10 
a = 8'd66; b = 8'd238;  #10 
a = 8'd66; b = 8'd239;  #10 
a = 8'd66; b = 8'd240;  #10 
a = 8'd66; b = 8'd241;  #10 
a = 8'd66; b = 8'd242;  #10 
a = 8'd66; b = 8'd243;  #10 
a = 8'd66; b = 8'd244;  #10 
a = 8'd66; b = 8'd245;  #10 
a = 8'd66; b = 8'd246;  #10 
a = 8'd66; b = 8'd247;  #10 
a = 8'd66; b = 8'd248;  #10 
a = 8'd66; b = 8'd249;  #10 
a = 8'd66; b = 8'd250;  #10 
a = 8'd66; b = 8'd251;  #10 
a = 8'd66; b = 8'd252;  #10 
a = 8'd66; b = 8'd253;  #10 
a = 8'd66; b = 8'd254;  #10 
a = 8'd66; b = 8'd255;  #10 
a = 8'd67; b = 8'd0;  #10 
a = 8'd67; b = 8'd1;  #10 
a = 8'd67; b = 8'd2;  #10 
a = 8'd67; b = 8'd3;  #10 
a = 8'd67; b = 8'd4;  #10 
a = 8'd67; b = 8'd5;  #10 
a = 8'd67; b = 8'd6;  #10 
a = 8'd67; b = 8'd7;  #10 
a = 8'd67; b = 8'd8;  #10 
a = 8'd67; b = 8'd9;  #10 
a = 8'd67; b = 8'd10;  #10 
a = 8'd67; b = 8'd11;  #10 
a = 8'd67; b = 8'd12;  #10 
a = 8'd67; b = 8'd13;  #10 
a = 8'd67; b = 8'd14;  #10 
a = 8'd67; b = 8'd15;  #10 
a = 8'd67; b = 8'd16;  #10 
a = 8'd67; b = 8'd17;  #10 
a = 8'd67; b = 8'd18;  #10 
a = 8'd67; b = 8'd19;  #10 
a = 8'd67; b = 8'd20;  #10 
a = 8'd67; b = 8'd21;  #10 
a = 8'd67; b = 8'd22;  #10 
a = 8'd67; b = 8'd23;  #10 
a = 8'd67; b = 8'd24;  #10 
a = 8'd67; b = 8'd25;  #10 
a = 8'd67; b = 8'd26;  #10 
a = 8'd67; b = 8'd27;  #10 
a = 8'd67; b = 8'd28;  #10 
a = 8'd67; b = 8'd29;  #10 
a = 8'd67; b = 8'd30;  #10 
a = 8'd67; b = 8'd31;  #10 
a = 8'd67; b = 8'd32;  #10 
a = 8'd67; b = 8'd33;  #10 
a = 8'd67; b = 8'd34;  #10 
a = 8'd67; b = 8'd35;  #10 
a = 8'd67; b = 8'd36;  #10 
a = 8'd67; b = 8'd37;  #10 
a = 8'd67; b = 8'd38;  #10 
a = 8'd67; b = 8'd39;  #10 
a = 8'd67; b = 8'd40;  #10 
a = 8'd67; b = 8'd41;  #10 
a = 8'd67; b = 8'd42;  #10 
a = 8'd67; b = 8'd43;  #10 
a = 8'd67; b = 8'd44;  #10 
a = 8'd67; b = 8'd45;  #10 
a = 8'd67; b = 8'd46;  #10 
a = 8'd67; b = 8'd47;  #10 
a = 8'd67; b = 8'd48;  #10 
a = 8'd67; b = 8'd49;  #10 
a = 8'd67; b = 8'd50;  #10 
a = 8'd67; b = 8'd51;  #10 
a = 8'd67; b = 8'd52;  #10 
a = 8'd67; b = 8'd53;  #10 
a = 8'd67; b = 8'd54;  #10 
a = 8'd67; b = 8'd55;  #10 
a = 8'd67; b = 8'd56;  #10 
a = 8'd67; b = 8'd57;  #10 
a = 8'd67; b = 8'd58;  #10 
a = 8'd67; b = 8'd59;  #10 
a = 8'd67; b = 8'd60;  #10 
a = 8'd67; b = 8'd61;  #10 
a = 8'd67; b = 8'd62;  #10 
a = 8'd67; b = 8'd63;  #10 
a = 8'd67; b = 8'd64;  #10 
a = 8'd67; b = 8'd65;  #10 
a = 8'd67; b = 8'd66;  #10 
a = 8'd67; b = 8'd67;  #10 
a = 8'd67; b = 8'd68;  #10 
a = 8'd67; b = 8'd69;  #10 
a = 8'd67; b = 8'd70;  #10 
a = 8'd67; b = 8'd71;  #10 
a = 8'd67; b = 8'd72;  #10 
a = 8'd67; b = 8'd73;  #10 
a = 8'd67; b = 8'd74;  #10 
a = 8'd67; b = 8'd75;  #10 
a = 8'd67; b = 8'd76;  #10 
a = 8'd67; b = 8'd77;  #10 
a = 8'd67; b = 8'd78;  #10 
a = 8'd67; b = 8'd79;  #10 
a = 8'd67; b = 8'd80;  #10 
a = 8'd67; b = 8'd81;  #10 
a = 8'd67; b = 8'd82;  #10 
a = 8'd67; b = 8'd83;  #10 
a = 8'd67; b = 8'd84;  #10 
a = 8'd67; b = 8'd85;  #10 
a = 8'd67; b = 8'd86;  #10 
a = 8'd67; b = 8'd87;  #10 
a = 8'd67; b = 8'd88;  #10 
a = 8'd67; b = 8'd89;  #10 
a = 8'd67; b = 8'd90;  #10 
a = 8'd67; b = 8'd91;  #10 
a = 8'd67; b = 8'd92;  #10 
a = 8'd67; b = 8'd93;  #10 
a = 8'd67; b = 8'd94;  #10 
a = 8'd67; b = 8'd95;  #10 
a = 8'd67; b = 8'd96;  #10 
a = 8'd67; b = 8'd97;  #10 
a = 8'd67; b = 8'd98;  #10 
a = 8'd67; b = 8'd99;  #10 
a = 8'd67; b = 8'd100;  #10 
a = 8'd67; b = 8'd101;  #10 
a = 8'd67; b = 8'd102;  #10 
a = 8'd67; b = 8'd103;  #10 
a = 8'd67; b = 8'd104;  #10 
a = 8'd67; b = 8'd105;  #10 
a = 8'd67; b = 8'd106;  #10 
a = 8'd67; b = 8'd107;  #10 
a = 8'd67; b = 8'd108;  #10 
a = 8'd67; b = 8'd109;  #10 
a = 8'd67; b = 8'd110;  #10 
a = 8'd67; b = 8'd111;  #10 
a = 8'd67; b = 8'd112;  #10 
a = 8'd67; b = 8'd113;  #10 
a = 8'd67; b = 8'd114;  #10 
a = 8'd67; b = 8'd115;  #10 
a = 8'd67; b = 8'd116;  #10 
a = 8'd67; b = 8'd117;  #10 
a = 8'd67; b = 8'd118;  #10 
a = 8'd67; b = 8'd119;  #10 
a = 8'd67; b = 8'd120;  #10 
a = 8'd67; b = 8'd121;  #10 
a = 8'd67; b = 8'd122;  #10 
a = 8'd67; b = 8'd123;  #10 
a = 8'd67; b = 8'd124;  #10 
a = 8'd67; b = 8'd125;  #10 
a = 8'd67; b = 8'd126;  #10 
a = 8'd67; b = 8'd127;  #10 
a = 8'd67; b = 8'd128;  #10 
a = 8'd67; b = 8'd129;  #10 
a = 8'd67; b = 8'd130;  #10 
a = 8'd67; b = 8'd131;  #10 
a = 8'd67; b = 8'd132;  #10 
a = 8'd67; b = 8'd133;  #10 
a = 8'd67; b = 8'd134;  #10 
a = 8'd67; b = 8'd135;  #10 
a = 8'd67; b = 8'd136;  #10 
a = 8'd67; b = 8'd137;  #10 
a = 8'd67; b = 8'd138;  #10 
a = 8'd67; b = 8'd139;  #10 
a = 8'd67; b = 8'd140;  #10 
a = 8'd67; b = 8'd141;  #10 
a = 8'd67; b = 8'd142;  #10 
a = 8'd67; b = 8'd143;  #10 
a = 8'd67; b = 8'd144;  #10 
a = 8'd67; b = 8'd145;  #10 
a = 8'd67; b = 8'd146;  #10 
a = 8'd67; b = 8'd147;  #10 
a = 8'd67; b = 8'd148;  #10 
a = 8'd67; b = 8'd149;  #10 
a = 8'd67; b = 8'd150;  #10 
a = 8'd67; b = 8'd151;  #10 
a = 8'd67; b = 8'd152;  #10 
a = 8'd67; b = 8'd153;  #10 
a = 8'd67; b = 8'd154;  #10 
a = 8'd67; b = 8'd155;  #10 
a = 8'd67; b = 8'd156;  #10 
a = 8'd67; b = 8'd157;  #10 
a = 8'd67; b = 8'd158;  #10 
a = 8'd67; b = 8'd159;  #10 
a = 8'd67; b = 8'd160;  #10 
a = 8'd67; b = 8'd161;  #10 
a = 8'd67; b = 8'd162;  #10 
a = 8'd67; b = 8'd163;  #10 
a = 8'd67; b = 8'd164;  #10 
a = 8'd67; b = 8'd165;  #10 
a = 8'd67; b = 8'd166;  #10 
a = 8'd67; b = 8'd167;  #10 
a = 8'd67; b = 8'd168;  #10 
a = 8'd67; b = 8'd169;  #10 
a = 8'd67; b = 8'd170;  #10 
a = 8'd67; b = 8'd171;  #10 
a = 8'd67; b = 8'd172;  #10 
a = 8'd67; b = 8'd173;  #10 
a = 8'd67; b = 8'd174;  #10 
a = 8'd67; b = 8'd175;  #10 
a = 8'd67; b = 8'd176;  #10 
a = 8'd67; b = 8'd177;  #10 
a = 8'd67; b = 8'd178;  #10 
a = 8'd67; b = 8'd179;  #10 
a = 8'd67; b = 8'd180;  #10 
a = 8'd67; b = 8'd181;  #10 
a = 8'd67; b = 8'd182;  #10 
a = 8'd67; b = 8'd183;  #10 
a = 8'd67; b = 8'd184;  #10 
a = 8'd67; b = 8'd185;  #10 
a = 8'd67; b = 8'd186;  #10 
a = 8'd67; b = 8'd187;  #10 
a = 8'd67; b = 8'd188;  #10 
a = 8'd67; b = 8'd189;  #10 
a = 8'd67; b = 8'd190;  #10 
a = 8'd67; b = 8'd191;  #10 
a = 8'd67; b = 8'd192;  #10 
a = 8'd67; b = 8'd193;  #10 
a = 8'd67; b = 8'd194;  #10 
a = 8'd67; b = 8'd195;  #10 
a = 8'd67; b = 8'd196;  #10 
a = 8'd67; b = 8'd197;  #10 
a = 8'd67; b = 8'd198;  #10 
a = 8'd67; b = 8'd199;  #10 
a = 8'd67; b = 8'd200;  #10 
a = 8'd67; b = 8'd201;  #10 
a = 8'd67; b = 8'd202;  #10 
a = 8'd67; b = 8'd203;  #10 
a = 8'd67; b = 8'd204;  #10 
a = 8'd67; b = 8'd205;  #10 
a = 8'd67; b = 8'd206;  #10 
a = 8'd67; b = 8'd207;  #10 
a = 8'd67; b = 8'd208;  #10 
a = 8'd67; b = 8'd209;  #10 
a = 8'd67; b = 8'd210;  #10 
a = 8'd67; b = 8'd211;  #10 
a = 8'd67; b = 8'd212;  #10 
a = 8'd67; b = 8'd213;  #10 
a = 8'd67; b = 8'd214;  #10 
a = 8'd67; b = 8'd215;  #10 
a = 8'd67; b = 8'd216;  #10 
a = 8'd67; b = 8'd217;  #10 
a = 8'd67; b = 8'd218;  #10 
a = 8'd67; b = 8'd219;  #10 
a = 8'd67; b = 8'd220;  #10 
a = 8'd67; b = 8'd221;  #10 
a = 8'd67; b = 8'd222;  #10 
a = 8'd67; b = 8'd223;  #10 
a = 8'd67; b = 8'd224;  #10 
a = 8'd67; b = 8'd225;  #10 
a = 8'd67; b = 8'd226;  #10 
a = 8'd67; b = 8'd227;  #10 
a = 8'd67; b = 8'd228;  #10 
a = 8'd67; b = 8'd229;  #10 
a = 8'd67; b = 8'd230;  #10 
a = 8'd67; b = 8'd231;  #10 
a = 8'd67; b = 8'd232;  #10 
a = 8'd67; b = 8'd233;  #10 
a = 8'd67; b = 8'd234;  #10 
a = 8'd67; b = 8'd235;  #10 
a = 8'd67; b = 8'd236;  #10 
a = 8'd67; b = 8'd237;  #10 
a = 8'd67; b = 8'd238;  #10 
a = 8'd67; b = 8'd239;  #10 
a = 8'd67; b = 8'd240;  #10 
a = 8'd67; b = 8'd241;  #10 
a = 8'd67; b = 8'd242;  #10 
a = 8'd67; b = 8'd243;  #10 
a = 8'd67; b = 8'd244;  #10 
a = 8'd67; b = 8'd245;  #10 
a = 8'd67; b = 8'd246;  #10 
a = 8'd67; b = 8'd247;  #10 
a = 8'd67; b = 8'd248;  #10 
a = 8'd67; b = 8'd249;  #10 
a = 8'd67; b = 8'd250;  #10 
a = 8'd67; b = 8'd251;  #10 
a = 8'd67; b = 8'd252;  #10 
a = 8'd67; b = 8'd253;  #10 
a = 8'd67; b = 8'd254;  #10 
a = 8'd67; b = 8'd255;  #10 
a = 8'd68; b = 8'd0;  #10 
a = 8'd68; b = 8'd1;  #10 
a = 8'd68; b = 8'd2;  #10 
a = 8'd68; b = 8'd3;  #10 
a = 8'd68; b = 8'd4;  #10 
a = 8'd68; b = 8'd5;  #10 
a = 8'd68; b = 8'd6;  #10 
a = 8'd68; b = 8'd7;  #10 
a = 8'd68; b = 8'd8;  #10 
a = 8'd68; b = 8'd9;  #10 
a = 8'd68; b = 8'd10;  #10 
a = 8'd68; b = 8'd11;  #10 
a = 8'd68; b = 8'd12;  #10 
a = 8'd68; b = 8'd13;  #10 
a = 8'd68; b = 8'd14;  #10 
a = 8'd68; b = 8'd15;  #10 
a = 8'd68; b = 8'd16;  #10 
a = 8'd68; b = 8'd17;  #10 
a = 8'd68; b = 8'd18;  #10 
a = 8'd68; b = 8'd19;  #10 
a = 8'd68; b = 8'd20;  #10 
a = 8'd68; b = 8'd21;  #10 
a = 8'd68; b = 8'd22;  #10 
a = 8'd68; b = 8'd23;  #10 
a = 8'd68; b = 8'd24;  #10 
a = 8'd68; b = 8'd25;  #10 
a = 8'd68; b = 8'd26;  #10 
a = 8'd68; b = 8'd27;  #10 
a = 8'd68; b = 8'd28;  #10 
a = 8'd68; b = 8'd29;  #10 
a = 8'd68; b = 8'd30;  #10 
a = 8'd68; b = 8'd31;  #10 
a = 8'd68; b = 8'd32;  #10 
a = 8'd68; b = 8'd33;  #10 
a = 8'd68; b = 8'd34;  #10 
a = 8'd68; b = 8'd35;  #10 
a = 8'd68; b = 8'd36;  #10 
a = 8'd68; b = 8'd37;  #10 
a = 8'd68; b = 8'd38;  #10 
a = 8'd68; b = 8'd39;  #10 
a = 8'd68; b = 8'd40;  #10 
a = 8'd68; b = 8'd41;  #10 
a = 8'd68; b = 8'd42;  #10 
a = 8'd68; b = 8'd43;  #10 
a = 8'd68; b = 8'd44;  #10 
a = 8'd68; b = 8'd45;  #10 
a = 8'd68; b = 8'd46;  #10 
a = 8'd68; b = 8'd47;  #10 
a = 8'd68; b = 8'd48;  #10 
a = 8'd68; b = 8'd49;  #10 
a = 8'd68; b = 8'd50;  #10 
a = 8'd68; b = 8'd51;  #10 
a = 8'd68; b = 8'd52;  #10 
a = 8'd68; b = 8'd53;  #10 
a = 8'd68; b = 8'd54;  #10 
a = 8'd68; b = 8'd55;  #10 
a = 8'd68; b = 8'd56;  #10 
a = 8'd68; b = 8'd57;  #10 
a = 8'd68; b = 8'd58;  #10 
a = 8'd68; b = 8'd59;  #10 
a = 8'd68; b = 8'd60;  #10 
a = 8'd68; b = 8'd61;  #10 
a = 8'd68; b = 8'd62;  #10 
a = 8'd68; b = 8'd63;  #10 
a = 8'd68; b = 8'd64;  #10 
a = 8'd68; b = 8'd65;  #10 
a = 8'd68; b = 8'd66;  #10 
a = 8'd68; b = 8'd67;  #10 
a = 8'd68; b = 8'd68;  #10 
a = 8'd68; b = 8'd69;  #10 
a = 8'd68; b = 8'd70;  #10 
a = 8'd68; b = 8'd71;  #10 
a = 8'd68; b = 8'd72;  #10 
a = 8'd68; b = 8'd73;  #10 
a = 8'd68; b = 8'd74;  #10 
a = 8'd68; b = 8'd75;  #10 
a = 8'd68; b = 8'd76;  #10 
a = 8'd68; b = 8'd77;  #10 
a = 8'd68; b = 8'd78;  #10 
a = 8'd68; b = 8'd79;  #10 
a = 8'd68; b = 8'd80;  #10 
a = 8'd68; b = 8'd81;  #10 
a = 8'd68; b = 8'd82;  #10 
a = 8'd68; b = 8'd83;  #10 
a = 8'd68; b = 8'd84;  #10 
a = 8'd68; b = 8'd85;  #10 
a = 8'd68; b = 8'd86;  #10 
a = 8'd68; b = 8'd87;  #10 
a = 8'd68; b = 8'd88;  #10 
a = 8'd68; b = 8'd89;  #10 
a = 8'd68; b = 8'd90;  #10 
a = 8'd68; b = 8'd91;  #10 
a = 8'd68; b = 8'd92;  #10 
a = 8'd68; b = 8'd93;  #10 
a = 8'd68; b = 8'd94;  #10 
a = 8'd68; b = 8'd95;  #10 
a = 8'd68; b = 8'd96;  #10 
a = 8'd68; b = 8'd97;  #10 
a = 8'd68; b = 8'd98;  #10 
a = 8'd68; b = 8'd99;  #10 
a = 8'd68; b = 8'd100;  #10 
a = 8'd68; b = 8'd101;  #10 
a = 8'd68; b = 8'd102;  #10 
a = 8'd68; b = 8'd103;  #10 
a = 8'd68; b = 8'd104;  #10 
a = 8'd68; b = 8'd105;  #10 
a = 8'd68; b = 8'd106;  #10 
a = 8'd68; b = 8'd107;  #10 
a = 8'd68; b = 8'd108;  #10 
a = 8'd68; b = 8'd109;  #10 
a = 8'd68; b = 8'd110;  #10 
a = 8'd68; b = 8'd111;  #10 
a = 8'd68; b = 8'd112;  #10 
a = 8'd68; b = 8'd113;  #10 
a = 8'd68; b = 8'd114;  #10 
a = 8'd68; b = 8'd115;  #10 
a = 8'd68; b = 8'd116;  #10 
a = 8'd68; b = 8'd117;  #10 
a = 8'd68; b = 8'd118;  #10 
a = 8'd68; b = 8'd119;  #10 
a = 8'd68; b = 8'd120;  #10 
a = 8'd68; b = 8'd121;  #10 
a = 8'd68; b = 8'd122;  #10 
a = 8'd68; b = 8'd123;  #10 
a = 8'd68; b = 8'd124;  #10 
a = 8'd68; b = 8'd125;  #10 
a = 8'd68; b = 8'd126;  #10 
a = 8'd68; b = 8'd127;  #10 
a = 8'd68; b = 8'd128;  #10 
a = 8'd68; b = 8'd129;  #10 
a = 8'd68; b = 8'd130;  #10 
a = 8'd68; b = 8'd131;  #10 
a = 8'd68; b = 8'd132;  #10 
a = 8'd68; b = 8'd133;  #10 
a = 8'd68; b = 8'd134;  #10 
a = 8'd68; b = 8'd135;  #10 
a = 8'd68; b = 8'd136;  #10 
a = 8'd68; b = 8'd137;  #10 
a = 8'd68; b = 8'd138;  #10 
a = 8'd68; b = 8'd139;  #10 
a = 8'd68; b = 8'd140;  #10 
a = 8'd68; b = 8'd141;  #10 
a = 8'd68; b = 8'd142;  #10 
a = 8'd68; b = 8'd143;  #10 
a = 8'd68; b = 8'd144;  #10 
a = 8'd68; b = 8'd145;  #10 
a = 8'd68; b = 8'd146;  #10 
a = 8'd68; b = 8'd147;  #10 
a = 8'd68; b = 8'd148;  #10 
a = 8'd68; b = 8'd149;  #10 
a = 8'd68; b = 8'd150;  #10 
a = 8'd68; b = 8'd151;  #10 
a = 8'd68; b = 8'd152;  #10 
a = 8'd68; b = 8'd153;  #10 
a = 8'd68; b = 8'd154;  #10 
a = 8'd68; b = 8'd155;  #10 
a = 8'd68; b = 8'd156;  #10 
a = 8'd68; b = 8'd157;  #10 
a = 8'd68; b = 8'd158;  #10 
a = 8'd68; b = 8'd159;  #10 
a = 8'd68; b = 8'd160;  #10 
a = 8'd68; b = 8'd161;  #10 
a = 8'd68; b = 8'd162;  #10 
a = 8'd68; b = 8'd163;  #10 
a = 8'd68; b = 8'd164;  #10 
a = 8'd68; b = 8'd165;  #10 
a = 8'd68; b = 8'd166;  #10 
a = 8'd68; b = 8'd167;  #10 
a = 8'd68; b = 8'd168;  #10 
a = 8'd68; b = 8'd169;  #10 
a = 8'd68; b = 8'd170;  #10 
a = 8'd68; b = 8'd171;  #10 
a = 8'd68; b = 8'd172;  #10 
a = 8'd68; b = 8'd173;  #10 
a = 8'd68; b = 8'd174;  #10 
a = 8'd68; b = 8'd175;  #10 
a = 8'd68; b = 8'd176;  #10 
a = 8'd68; b = 8'd177;  #10 
a = 8'd68; b = 8'd178;  #10 
a = 8'd68; b = 8'd179;  #10 
a = 8'd68; b = 8'd180;  #10 
a = 8'd68; b = 8'd181;  #10 
a = 8'd68; b = 8'd182;  #10 
a = 8'd68; b = 8'd183;  #10 
a = 8'd68; b = 8'd184;  #10 
a = 8'd68; b = 8'd185;  #10 
a = 8'd68; b = 8'd186;  #10 
a = 8'd68; b = 8'd187;  #10 
a = 8'd68; b = 8'd188;  #10 
a = 8'd68; b = 8'd189;  #10 
a = 8'd68; b = 8'd190;  #10 
a = 8'd68; b = 8'd191;  #10 
a = 8'd68; b = 8'd192;  #10 
a = 8'd68; b = 8'd193;  #10 
a = 8'd68; b = 8'd194;  #10 
a = 8'd68; b = 8'd195;  #10 
a = 8'd68; b = 8'd196;  #10 
a = 8'd68; b = 8'd197;  #10 
a = 8'd68; b = 8'd198;  #10 
a = 8'd68; b = 8'd199;  #10 
a = 8'd68; b = 8'd200;  #10 
a = 8'd68; b = 8'd201;  #10 
a = 8'd68; b = 8'd202;  #10 
a = 8'd68; b = 8'd203;  #10 
a = 8'd68; b = 8'd204;  #10 
a = 8'd68; b = 8'd205;  #10 
a = 8'd68; b = 8'd206;  #10 
a = 8'd68; b = 8'd207;  #10 
a = 8'd68; b = 8'd208;  #10 
a = 8'd68; b = 8'd209;  #10 
a = 8'd68; b = 8'd210;  #10 
a = 8'd68; b = 8'd211;  #10 
a = 8'd68; b = 8'd212;  #10 
a = 8'd68; b = 8'd213;  #10 
a = 8'd68; b = 8'd214;  #10 
a = 8'd68; b = 8'd215;  #10 
a = 8'd68; b = 8'd216;  #10 
a = 8'd68; b = 8'd217;  #10 
a = 8'd68; b = 8'd218;  #10 
a = 8'd68; b = 8'd219;  #10 
a = 8'd68; b = 8'd220;  #10 
a = 8'd68; b = 8'd221;  #10 
a = 8'd68; b = 8'd222;  #10 
a = 8'd68; b = 8'd223;  #10 
a = 8'd68; b = 8'd224;  #10 
a = 8'd68; b = 8'd225;  #10 
a = 8'd68; b = 8'd226;  #10 
a = 8'd68; b = 8'd227;  #10 
a = 8'd68; b = 8'd228;  #10 
a = 8'd68; b = 8'd229;  #10 
a = 8'd68; b = 8'd230;  #10 
a = 8'd68; b = 8'd231;  #10 
a = 8'd68; b = 8'd232;  #10 
a = 8'd68; b = 8'd233;  #10 
a = 8'd68; b = 8'd234;  #10 
a = 8'd68; b = 8'd235;  #10 
a = 8'd68; b = 8'd236;  #10 
a = 8'd68; b = 8'd237;  #10 
a = 8'd68; b = 8'd238;  #10 
a = 8'd68; b = 8'd239;  #10 
a = 8'd68; b = 8'd240;  #10 
a = 8'd68; b = 8'd241;  #10 
a = 8'd68; b = 8'd242;  #10 
a = 8'd68; b = 8'd243;  #10 
a = 8'd68; b = 8'd244;  #10 
a = 8'd68; b = 8'd245;  #10 
a = 8'd68; b = 8'd246;  #10 
a = 8'd68; b = 8'd247;  #10 
a = 8'd68; b = 8'd248;  #10 
a = 8'd68; b = 8'd249;  #10 
a = 8'd68; b = 8'd250;  #10 
a = 8'd68; b = 8'd251;  #10 
a = 8'd68; b = 8'd252;  #10 
a = 8'd68; b = 8'd253;  #10 
a = 8'd68; b = 8'd254;  #10 
a = 8'd68; b = 8'd255;  #10 
a = 8'd69; b = 8'd0;  #10 
a = 8'd69; b = 8'd1;  #10 
a = 8'd69; b = 8'd2;  #10 
a = 8'd69; b = 8'd3;  #10 
a = 8'd69; b = 8'd4;  #10 
a = 8'd69; b = 8'd5;  #10 
a = 8'd69; b = 8'd6;  #10 
a = 8'd69; b = 8'd7;  #10 
a = 8'd69; b = 8'd8;  #10 
a = 8'd69; b = 8'd9;  #10 
a = 8'd69; b = 8'd10;  #10 
a = 8'd69; b = 8'd11;  #10 
a = 8'd69; b = 8'd12;  #10 
a = 8'd69; b = 8'd13;  #10 
a = 8'd69; b = 8'd14;  #10 
a = 8'd69; b = 8'd15;  #10 
a = 8'd69; b = 8'd16;  #10 
a = 8'd69; b = 8'd17;  #10 
a = 8'd69; b = 8'd18;  #10 
a = 8'd69; b = 8'd19;  #10 
a = 8'd69; b = 8'd20;  #10 
a = 8'd69; b = 8'd21;  #10 
a = 8'd69; b = 8'd22;  #10 
a = 8'd69; b = 8'd23;  #10 
a = 8'd69; b = 8'd24;  #10 
a = 8'd69; b = 8'd25;  #10 
a = 8'd69; b = 8'd26;  #10 
a = 8'd69; b = 8'd27;  #10 
a = 8'd69; b = 8'd28;  #10 
a = 8'd69; b = 8'd29;  #10 
a = 8'd69; b = 8'd30;  #10 
a = 8'd69; b = 8'd31;  #10 
a = 8'd69; b = 8'd32;  #10 
a = 8'd69; b = 8'd33;  #10 
a = 8'd69; b = 8'd34;  #10 
a = 8'd69; b = 8'd35;  #10 
a = 8'd69; b = 8'd36;  #10 
a = 8'd69; b = 8'd37;  #10 
a = 8'd69; b = 8'd38;  #10 
a = 8'd69; b = 8'd39;  #10 
a = 8'd69; b = 8'd40;  #10 
a = 8'd69; b = 8'd41;  #10 
a = 8'd69; b = 8'd42;  #10 
a = 8'd69; b = 8'd43;  #10 
a = 8'd69; b = 8'd44;  #10 
a = 8'd69; b = 8'd45;  #10 
a = 8'd69; b = 8'd46;  #10 
a = 8'd69; b = 8'd47;  #10 
a = 8'd69; b = 8'd48;  #10 
a = 8'd69; b = 8'd49;  #10 
a = 8'd69; b = 8'd50;  #10 
a = 8'd69; b = 8'd51;  #10 
a = 8'd69; b = 8'd52;  #10 
a = 8'd69; b = 8'd53;  #10 
a = 8'd69; b = 8'd54;  #10 
a = 8'd69; b = 8'd55;  #10 
a = 8'd69; b = 8'd56;  #10 
a = 8'd69; b = 8'd57;  #10 
a = 8'd69; b = 8'd58;  #10 
a = 8'd69; b = 8'd59;  #10 
a = 8'd69; b = 8'd60;  #10 
a = 8'd69; b = 8'd61;  #10 
a = 8'd69; b = 8'd62;  #10 
a = 8'd69; b = 8'd63;  #10 
a = 8'd69; b = 8'd64;  #10 
a = 8'd69; b = 8'd65;  #10 
a = 8'd69; b = 8'd66;  #10 
a = 8'd69; b = 8'd67;  #10 
a = 8'd69; b = 8'd68;  #10 
a = 8'd69; b = 8'd69;  #10 
a = 8'd69; b = 8'd70;  #10 
a = 8'd69; b = 8'd71;  #10 
a = 8'd69; b = 8'd72;  #10 
a = 8'd69; b = 8'd73;  #10 
a = 8'd69; b = 8'd74;  #10 
a = 8'd69; b = 8'd75;  #10 
a = 8'd69; b = 8'd76;  #10 
a = 8'd69; b = 8'd77;  #10 
a = 8'd69; b = 8'd78;  #10 
a = 8'd69; b = 8'd79;  #10 
a = 8'd69; b = 8'd80;  #10 
a = 8'd69; b = 8'd81;  #10 
a = 8'd69; b = 8'd82;  #10 
a = 8'd69; b = 8'd83;  #10 
a = 8'd69; b = 8'd84;  #10 
a = 8'd69; b = 8'd85;  #10 
a = 8'd69; b = 8'd86;  #10 
a = 8'd69; b = 8'd87;  #10 
a = 8'd69; b = 8'd88;  #10 
a = 8'd69; b = 8'd89;  #10 
a = 8'd69; b = 8'd90;  #10 
a = 8'd69; b = 8'd91;  #10 
a = 8'd69; b = 8'd92;  #10 
a = 8'd69; b = 8'd93;  #10 
a = 8'd69; b = 8'd94;  #10 
a = 8'd69; b = 8'd95;  #10 
a = 8'd69; b = 8'd96;  #10 
a = 8'd69; b = 8'd97;  #10 
a = 8'd69; b = 8'd98;  #10 
a = 8'd69; b = 8'd99;  #10 
a = 8'd69; b = 8'd100;  #10 
a = 8'd69; b = 8'd101;  #10 
a = 8'd69; b = 8'd102;  #10 
a = 8'd69; b = 8'd103;  #10 
a = 8'd69; b = 8'd104;  #10 
a = 8'd69; b = 8'd105;  #10 
a = 8'd69; b = 8'd106;  #10 
a = 8'd69; b = 8'd107;  #10 
a = 8'd69; b = 8'd108;  #10 
a = 8'd69; b = 8'd109;  #10 
a = 8'd69; b = 8'd110;  #10 
a = 8'd69; b = 8'd111;  #10 
a = 8'd69; b = 8'd112;  #10 
a = 8'd69; b = 8'd113;  #10 
a = 8'd69; b = 8'd114;  #10 
a = 8'd69; b = 8'd115;  #10 
a = 8'd69; b = 8'd116;  #10 
a = 8'd69; b = 8'd117;  #10 
a = 8'd69; b = 8'd118;  #10 
a = 8'd69; b = 8'd119;  #10 
a = 8'd69; b = 8'd120;  #10 
a = 8'd69; b = 8'd121;  #10 
a = 8'd69; b = 8'd122;  #10 
a = 8'd69; b = 8'd123;  #10 
a = 8'd69; b = 8'd124;  #10 
a = 8'd69; b = 8'd125;  #10 
a = 8'd69; b = 8'd126;  #10 
a = 8'd69; b = 8'd127;  #10 
a = 8'd69; b = 8'd128;  #10 
a = 8'd69; b = 8'd129;  #10 
a = 8'd69; b = 8'd130;  #10 
a = 8'd69; b = 8'd131;  #10 
a = 8'd69; b = 8'd132;  #10 
a = 8'd69; b = 8'd133;  #10 
a = 8'd69; b = 8'd134;  #10 
a = 8'd69; b = 8'd135;  #10 
a = 8'd69; b = 8'd136;  #10 
a = 8'd69; b = 8'd137;  #10 
a = 8'd69; b = 8'd138;  #10 
a = 8'd69; b = 8'd139;  #10 
a = 8'd69; b = 8'd140;  #10 
a = 8'd69; b = 8'd141;  #10 
a = 8'd69; b = 8'd142;  #10 
a = 8'd69; b = 8'd143;  #10 
a = 8'd69; b = 8'd144;  #10 
a = 8'd69; b = 8'd145;  #10 
a = 8'd69; b = 8'd146;  #10 
a = 8'd69; b = 8'd147;  #10 
a = 8'd69; b = 8'd148;  #10 
a = 8'd69; b = 8'd149;  #10 
a = 8'd69; b = 8'd150;  #10 
a = 8'd69; b = 8'd151;  #10 
a = 8'd69; b = 8'd152;  #10 
a = 8'd69; b = 8'd153;  #10 
a = 8'd69; b = 8'd154;  #10 
a = 8'd69; b = 8'd155;  #10 
a = 8'd69; b = 8'd156;  #10 
a = 8'd69; b = 8'd157;  #10 
a = 8'd69; b = 8'd158;  #10 
a = 8'd69; b = 8'd159;  #10 
a = 8'd69; b = 8'd160;  #10 
a = 8'd69; b = 8'd161;  #10 
a = 8'd69; b = 8'd162;  #10 
a = 8'd69; b = 8'd163;  #10 
a = 8'd69; b = 8'd164;  #10 
a = 8'd69; b = 8'd165;  #10 
a = 8'd69; b = 8'd166;  #10 
a = 8'd69; b = 8'd167;  #10 
a = 8'd69; b = 8'd168;  #10 
a = 8'd69; b = 8'd169;  #10 
a = 8'd69; b = 8'd170;  #10 
a = 8'd69; b = 8'd171;  #10 
a = 8'd69; b = 8'd172;  #10 
a = 8'd69; b = 8'd173;  #10 
a = 8'd69; b = 8'd174;  #10 
a = 8'd69; b = 8'd175;  #10 
a = 8'd69; b = 8'd176;  #10 
a = 8'd69; b = 8'd177;  #10 
a = 8'd69; b = 8'd178;  #10 
a = 8'd69; b = 8'd179;  #10 
a = 8'd69; b = 8'd180;  #10 
a = 8'd69; b = 8'd181;  #10 
a = 8'd69; b = 8'd182;  #10 
a = 8'd69; b = 8'd183;  #10 
a = 8'd69; b = 8'd184;  #10 
a = 8'd69; b = 8'd185;  #10 
a = 8'd69; b = 8'd186;  #10 
a = 8'd69; b = 8'd187;  #10 
a = 8'd69; b = 8'd188;  #10 
a = 8'd69; b = 8'd189;  #10 
a = 8'd69; b = 8'd190;  #10 
a = 8'd69; b = 8'd191;  #10 
a = 8'd69; b = 8'd192;  #10 
a = 8'd69; b = 8'd193;  #10 
a = 8'd69; b = 8'd194;  #10 
a = 8'd69; b = 8'd195;  #10 
a = 8'd69; b = 8'd196;  #10 
a = 8'd69; b = 8'd197;  #10 
a = 8'd69; b = 8'd198;  #10 
a = 8'd69; b = 8'd199;  #10 
a = 8'd69; b = 8'd200;  #10 
a = 8'd69; b = 8'd201;  #10 
a = 8'd69; b = 8'd202;  #10 
a = 8'd69; b = 8'd203;  #10 
a = 8'd69; b = 8'd204;  #10 
a = 8'd69; b = 8'd205;  #10 
a = 8'd69; b = 8'd206;  #10 
a = 8'd69; b = 8'd207;  #10 
a = 8'd69; b = 8'd208;  #10 
a = 8'd69; b = 8'd209;  #10 
a = 8'd69; b = 8'd210;  #10 
a = 8'd69; b = 8'd211;  #10 
a = 8'd69; b = 8'd212;  #10 
a = 8'd69; b = 8'd213;  #10 
a = 8'd69; b = 8'd214;  #10 
a = 8'd69; b = 8'd215;  #10 
a = 8'd69; b = 8'd216;  #10 
a = 8'd69; b = 8'd217;  #10 
a = 8'd69; b = 8'd218;  #10 
a = 8'd69; b = 8'd219;  #10 
a = 8'd69; b = 8'd220;  #10 
a = 8'd69; b = 8'd221;  #10 
a = 8'd69; b = 8'd222;  #10 
a = 8'd69; b = 8'd223;  #10 
a = 8'd69; b = 8'd224;  #10 
a = 8'd69; b = 8'd225;  #10 
a = 8'd69; b = 8'd226;  #10 
a = 8'd69; b = 8'd227;  #10 
a = 8'd69; b = 8'd228;  #10 
a = 8'd69; b = 8'd229;  #10 
a = 8'd69; b = 8'd230;  #10 
a = 8'd69; b = 8'd231;  #10 
a = 8'd69; b = 8'd232;  #10 
a = 8'd69; b = 8'd233;  #10 
a = 8'd69; b = 8'd234;  #10 
a = 8'd69; b = 8'd235;  #10 
a = 8'd69; b = 8'd236;  #10 
a = 8'd69; b = 8'd237;  #10 
a = 8'd69; b = 8'd238;  #10 
a = 8'd69; b = 8'd239;  #10 
a = 8'd69; b = 8'd240;  #10 
a = 8'd69; b = 8'd241;  #10 
a = 8'd69; b = 8'd242;  #10 
a = 8'd69; b = 8'd243;  #10 
a = 8'd69; b = 8'd244;  #10 
a = 8'd69; b = 8'd245;  #10 
a = 8'd69; b = 8'd246;  #10 
a = 8'd69; b = 8'd247;  #10 
a = 8'd69; b = 8'd248;  #10 
a = 8'd69; b = 8'd249;  #10 
a = 8'd69; b = 8'd250;  #10 
a = 8'd69; b = 8'd251;  #10 
a = 8'd69; b = 8'd252;  #10 
a = 8'd69; b = 8'd253;  #10 
a = 8'd69; b = 8'd254;  #10 
a = 8'd69; b = 8'd255;  #10 
a = 8'd70; b = 8'd0;  #10 
a = 8'd70; b = 8'd1;  #10 
a = 8'd70; b = 8'd2;  #10 
a = 8'd70; b = 8'd3;  #10 
a = 8'd70; b = 8'd4;  #10 
a = 8'd70; b = 8'd5;  #10 
a = 8'd70; b = 8'd6;  #10 
a = 8'd70; b = 8'd7;  #10 
a = 8'd70; b = 8'd8;  #10 
a = 8'd70; b = 8'd9;  #10 
a = 8'd70; b = 8'd10;  #10 
a = 8'd70; b = 8'd11;  #10 
a = 8'd70; b = 8'd12;  #10 
a = 8'd70; b = 8'd13;  #10 
a = 8'd70; b = 8'd14;  #10 
a = 8'd70; b = 8'd15;  #10 
a = 8'd70; b = 8'd16;  #10 
a = 8'd70; b = 8'd17;  #10 
a = 8'd70; b = 8'd18;  #10 
a = 8'd70; b = 8'd19;  #10 
a = 8'd70; b = 8'd20;  #10 
a = 8'd70; b = 8'd21;  #10 
a = 8'd70; b = 8'd22;  #10 
a = 8'd70; b = 8'd23;  #10 
a = 8'd70; b = 8'd24;  #10 
a = 8'd70; b = 8'd25;  #10 
a = 8'd70; b = 8'd26;  #10 
a = 8'd70; b = 8'd27;  #10 
a = 8'd70; b = 8'd28;  #10 
a = 8'd70; b = 8'd29;  #10 
a = 8'd70; b = 8'd30;  #10 
a = 8'd70; b = 8'd31;  #10 
a = 8'd70; b = 8'd32;  #10 
a = 8'd70; b = 8'd33;  #10 
a = 8'd70; b = 8'd34;  #10 
a = 8'd70; b = 8'd35;  #10 
a = 8'd70; b = 8'd36;  #10 
a = 8'd70; b = 8'd37;  #10 
a = 8'd70; b = 8'd38;  #10 
a = 8'd70; b = 8'd39;  #10 
a = 8'd70; b = 8'd40;  #10 
a = 8'd70; b = 8'd41;  #10 
a = 8'd70; b = 8'd42;  #10 
a = 8'd70; b = 8'd43;  #10 
a = 8'd70; b = 8'd44;  #10 
a = 8'd70; b = 8'd45;  #10 
a = 8'd70; b = 8'd46;  #10 
a = 8'd70; b = 8'd47;  #10 
a = 8'd70; b = 8'd48;  #10 
a = 8'd70; b = 8'd49;  #10 
a = 8'd70; b = 8'd50;  #10 
a = 8'd70; b = 8'd51;  #10 
a = 8'd70; b = 8'd52;  #10 
a = 8'd70; b = 8'd53;  #10 
a = 8'd70; b = 8'd54;  #10 
a = 8'd70; b = 8'd55;  #10 
a = 8'd70; b = 8'd56;  #10 
a = 8'd70; b = 8'd57;  #10 
a = 8'd70; b = 8'd58;  #10 
a = 8'd70; b = 8'd59;  #10 
a = 8'd70; b = 8'd60;  #10 
a = 8'd70; b = 8'd61;  #10 
a = 8'd70; b = 8'd62;  #10 
a = 8'd70; b = 8'd63;  #10 
a = 8'd70; b = 8'd64;  #10 
a = 8'd70; b = 8'd65;  #10 
a = 8'd70; b = 8'd66;  #10 
a = 8'd70; b = 8'd67;  #10 
a = 8'd70; b = 8'd68;  #10 
a = 8'd70; b = 8'd69;  #10 
a = 8'd70; b = 8'd70;  #10 
a = 8'd70; b = 8'd71;  #10 
a = 8'd70; b = 8'd72;  #10 
a = 8'd70; b = 8'd73;  #10 
a = 8'd70; b = 8'd74;  #10 
a = 8'd70; b = 8'd75;  #10 
a = 8'd70; b = 8'd76;  #10 
a = 8'd70; b = 8'd77;  #10 
a = 8'd70; b = 8'd78;  #10 
a = 8'd70; b = 8'd79;  #10 
a = 8'd70; b = 8'd80;  #10 
a = 8'd70; b = 8'd81;  #10 
a = 8'd70; b = 8'd82;  #10 
a = 8'd70; b = 8'd83;  #10 
a = 8'd70; b = 8'd84;  #10 
a = 8'd70; b = 8'd85;  #10 
a = 8'd70; b = 8'd86;  #10 
a = 8'd70; b = 8'd87;  #10 
a = 8'd70; b = 8'd88;  #10 
a = 8'd70; b = 8'd89;  #10 
a = 8'd70; b = 8'd90;  #10 
a = 8'd70; b = 8'd91;  #10 
a = 8'd70; b = 8'd92;  #10 
a = 8'd70; b = 8'd93;  #10 
a = 8'd70; b = 8'd94;  #10 
a = 8'd70; b = 8'd95;  #10 
a = 8'd70; b = 8'd96;  #10 
a = 8'd70; b = 8'd97;  #10 
a = 8'd70; b = 8'd98;  #10 
a = 8'd70; b = 8'd99;  #10 
a = 8'd70; b = 8'd100;  #10 
a = 8'd70; b = 8'd101;  #10 
a = 8'd70; b = 8'd102;  #10 
a = 8'd70; b = 8'd103;  #10 
a = 8'd70; b = 8'd104;  #10 
a = 8'd70; b = 8'd105;  #10 
a = 8'd70; b = 8'd106;  #10 
a = 8'd70; b = 8'd107;  #10 
a = 8'd70; b = 8'd108;  #10 
a = 8'd70; b = 8'd109;  #10 
a = 8'd70; b = 8'd110;  #10 
a = 8'd70; b = 8'd111;  #10 
a = 8'd70; b = 8'd112;  #10 
a = 8'd70; b = 8'd113;  #10 
a = 8'd70; b = 8'd114;  #10 
a = 8'd70; b = 8'd115;  #10 
a = 8'd70; b = 8'd116;  #10 
a = 8'd70; b = 8'd117;  #10 
a = 8'd70; b = 8'd118;  #10 
a = 8'd70; b = 8'd119;  #10 
a = 8'd70; b = 8'd120;  #10 
a = 8'd70; b = 8'd121;  #10 
a = 8'd70; b = 8'd122;  #10 
a = 8'd70; b = 8'd123;  #10 
a = 8'd70; b = 8'd124;  #10 
a = 8'd70; b = 8'd125;  #10 
a = 8'd70; b = 8'd126;  #10 
a = 8'd70; b = 8'd127;  #10 
a = 8'd70; b = 8'd128;  #10 
a = 8'd70; b = 8'd129;  #10 
a = 8'd70; b = 8'd130;  #10 
a = 8'd70; b = 8'd131;  #10 
a = 8'd70; b = 8'd132;  #10 
a = 8'd70; b = 8'd133;  #10 
a = 8'd70; b = 8'd134;  #10 
a = 8'd70; b = 8'd135;  #10 
a = 8'd70; b = 8'd136;  #10 
a = 8'd70; b = 8'd137;  #10 
a = 8'd70; b = 8'd138;  #10 
a = 8'd70; b = 8'd139;  #10 
a = 8'd70; b = 8'd140;  #10 
a = 8'd70; b = 8'd141;  #10 
a = 8'd70; b = 8'd142;  #10 
a = 8'd70; b = 8'd143;  #10 
a = 8'd70; b = 8'd144;  #10 
a = 8'd70; b = 8'd145;  #10 
a = 8'd70; b = 8'd146;  #10 
a = 8'd70; b = 8'd147;  #10 
a = 8'd70; b = 8'd148;  #10 
a = 8'd70; b = 8'd149;  #10 
a = 8'd70; b = 8'd150;  #10 
a = 8'd70; b = 8'd151;  #10 
a = 8'd70; b = 8'd152;  #10 
a = 8'd70; b = 8'd153;  #10 
a = 8'd70; b = 8'd154;  #10 
a = 8'd70; b = 8'd155;  #10 
a = 8'd70; b = 8'd156;  #10 
a = 8'd70; b = 8'd157;  #10 
a = 8'd70; b = 8'd158;  #10 
a = 8'd70; b = 8'd159;  #10 
a = 8'd70; b = 8'd160;  #10 
a = 8'd70; b = 8'd161;  #10 
a = 8'd70; b = 8'd162;  #10 
a = 8'd70; b = 8'd163;  #10 
a = 8'd70; b = 8'd164;  #10 
a = 8'd70; b = 8'd165;  #10 
a = 8'd70; b = 8'd166;  #10 
a = 8'd70; b = 8'd167;  #10 
a = 8'd70; b = 8'd168;  #10 
a = 8'd70; b = 8'd169;  #10 
a = 8'd70; b = 8'd170;  #10 
a = 8'd70; b = 8'd171;  #10 
a = 8'd70; b = 8'd172;  #10 
a = 8'd70; b = 8'd173;  #10 
a = 8'd70; b = 8'd174;  #10 
a = 8'd70; b = 8'd175;  #10 
a = 8'd70; b = 8'd176;  #10 
a = 8'd70; b = 8'd177;  #10 
a = 8'd70; b = 8'd178;  #10 
a = 8'd70; b = 8'd179;  #10 
a = 8'd70; b = 8'd180;  #10 
a = 8'd70; b = 8'd181;  #10 
a = 8'd70; b = 8'd182;  #10 
a = 8'd70; b = 8'd183;  #10 
a = 8'd70; b = 8'd184;  #10 
a = 8'd70; b = 8'd185;  #10 
a = 8'd70; b = 8'd186;  #10 
a = 8'd70; b = 8'd187;  #10 
a = 8'd70; b = 8'd188;  #10 
a = 8'd70; b = 8'd189;  #10 
a = 8'd70; b = 8'd190;  #10 
a = 8'd70; b = 8'd191;  #10 
a = 8'd70; b = 8'd192;  #10 
a = 8'd70; b = 8'd193;  #10 
a = 8'd70; b = 8'd194;  #10 
a = 8'd70; b = 8'd195;  #10 
a = 8'd70; b = 8'd196;  #10 
a = 8'd70; b = 8'd197;  #10 
a = 8'd70; b = 8'd198;  #10 
a = 8'd70; b = 8'd199;  #10 
a = 8'd70; b = 8'd200;  #10 
a = 8'd70; b = 8'd201;  #10 
a = 8'd70; b = 8'd202;  #10 
a = 8'd70; b = 8'd203;  #10 
a = 8'd70; b = 8'd204;  #10 
a = 8'd70; b = 8'd205;  #10 
a = 8'd70; b = 8'd206;  #10 
a = 8'd70; b = 8'd207;  #10 
a = 8'd70; b = 8'd208;  #10 
a = 8'd70; b = 8'd209;  #10 
a = 8'd70; b = 8'd210;  #10 
a = 8'd70; b = 8'd211;  #10 
a = 8'd70; b = 8'd212;  #10 
a = 8'd70; b = 8'd213;  #10 
a = 8'd70; b = 8'd214;  #10 
a = 8'd70; b = 8'd215;  #10 
a = 8'd70; b = 8'd216;  #10 
a = 8'd70; b = 8'd217;  #10 
a = 8'd70; b = 8'd218;  #10 
a = 8'd70; b = 8'd219;  #10 
a = 8'd70; b = 8'd220;  #10 
a = 8'd70; b = 8'd221;  #10 
a = 8'd70; b = 8'd222;  #10 
a = 8'd70; b = 8'd223;  #10 
a = 8'd70; b = 8'd224;  #10 
a = 8'd70; b = 8'd225;  #10 
a = 8'd70; b = 8'd226;  #10 
a = 8'd70; b = 8'd227;  #10 
a = 8'd70; b = 8'd228;  #10 
a = 8'd70; b = 8'd229;  #10 
a = 8'd70; b = 8'd230;  #10 
a = 8'd70; b = 8'd231;  #10 
a = 8'd70; b = 8'd232;  #10 
a = 8'd70; b = 8'd233;  #10 
a = 8'd70; b = 8'd234;  #10 
a = 8'd70; b = 8'd235;  #10 
a = 8'd70; b = 8'd236;  #10 
a = 8'd70; b = 8'd237;  #10 
a = 8'd70; b = 8'd238;  #10 
a = 8'd70; b = 8'd239;  #10 
a = 8'd70; b = 8'd240;  #10 
a = 8'd70; b = 8'd241;  #10 
a = 8'd70; b = 8'd242;  #10 
a = 8'd70; b = 8'd243;  #10 
a = 8'd70; b = 8'd244;  #10 
a = 8'd70; b = 8'd245;  #10 
a = 8'd70; b = 8'd246;  #10 
a = 8'd70; b = 8'd247;  #10 
a = 8'd70; b = 8'd248;  #10 
a = 8'd70; b = 8'd249;  #10 
a = 8'd70; b = 8'd250;  #10 
a = 8'd70; b = 8'd251;  #10 
a = 8'd70; b = 8'd252;  #10 
a = 8'd70; b = 8'd253;  #10 
a = 8'd70; b = 8'd254;  #10 
a = 8'd70; b = 8'd255;  #10 
a = 8'd71; b = 8'd0;  #10 
a = 8'd71; b = 8'd1;  #10 
a = 8'd71; b = 8'd2;  #10 
a = 8'd71; b = 8'd3;  #10 
a = 8'd71; b = 8'd4;  #10 
a = 8'd71; b = 8'd5;  #10 
a = 8'd71; b = 8'd6;  #10 
a = 8'd71; b = 8'd7;  #10 
a = 8'd71; b = 8'd8;  #10 
a = 8'd71; b = 8'd9;  #10 
a = 8'd71; b = 8'd10;  #10 
a = 8'd71; b = 8'd11;  #10 
a = 8'd71; b = 8'd12;  #10 
a = 8'd71; b = 8'd13;  #10 
a = 8'd71; b = 8'd14;  #10 
a = 8'd71; b = 8'd15;  #10 
a = 8'd71; b = 8'd16;  #10 
a = 8'd71; b = 8'd17;  #10 
a = 8'd71; b = 8'd18;  #10 
a = 8'd71; b = 8'd19;  #10 
a = 8'd71; b = 8'd20;  #10 
a = 8'd71; b = 8'd21;  #10 
a = 8'd71; b = 8'd22;  #10 
a = 8'd71; b = 8'd23;  #10 
a = 8'd71; b = 8'd24;  #10 
a = 8'd71; b = 8'd25;  #10 
a = 8'd71; b = 8'd26;  #10 
a = 8'd71; b = 8'd27;  #10 
a = 8'd71; b = 8'd28;  #10 
a = 8'd71; b = 8'd29;  #10 
a = 8'd71; b = 8'd30;  #10 
a = 8'd71; b = 8'd31;  #10 
a = 8'd71; b = 8'd32;  #10 
a = 8'd71; b = 8'd33;  #10 
a = 8'd71; b = 8'd34;  #10 
a = 8'd71; b = 8'd35;  #10 
a = 8'd71; b = 8'd36;  #10 
a = 8'd71; b = 8'd37;  #10 
a = 8'd71; b = 8'd38;  #10 
a = 8'd71; b = 8'd39;  #10 
a = 8'd71; b = 8'd40;  #10 
a = 8'd71; b = 8'd41;  #10 
a = 8'd71; b = 8'd42;  #10 
a = 8'd71; b = 8'd43;  #10 
a = 8'd71; b = 8'd44;  #10 
a = 8'd71; b = 8'd45;  #10 
a = 8'd71; b = 8'd46;  #10 
a = 8'd71; b = 8'd47;  #10 
a = 8'd71; b = 8'd48;  #10 
a = 8'd71; b = 8'd49;  #10 
a = 8'd71; b = 8'd50;  #10 
a = 8'd71; b = 8'd51;  #10 
a = 8'd71; b = 8'd52;  #10 
a = 8'd71; b = 8'd53;  #10 
a = 8'd71; b = 8'd54;  #10 
a = 8'd71; b = 8'd55;  #10 
a = 8'd71; b = 8'd56;  #10 
a = 8'd71; b = 8'd57;  #10 
a = 8'd71; b = 8'd58;  #10 
a = 8'd71; b = 8'd59;  #10 
a = 8'd71; b = 8'd60;  #10 
a = 8'd71; b = 8'd61;  #10 
a = 8'd71; b = 8'd62;  #10 
a = 8'd71; b = 8'd63;  #10 
a = 8'd71; b = 8'd64;  #10 
a = 8'd71; b = 8'd65;  #10 
a = 8'd71; b = 8'd66;  #10 
a = 8'd71; b = 8'd67;  #10 
a = 8'd71; b = 8'd68;  #10 
a = 8'd71; b = 8'd69;  #10 
a = 8'd71; b = 8'd70;  #10 
a = 8'd71; b = 8'd71;  #10 
a = 8'd71; b = 8'd72;  #10 
a = 8'd71; b = 8'd73;  #10 
a = 8'd71; b = 8'd74;  #10 
a = 8'd71; b = 8'd75;  #10 
a = 8'd71; b = 8'd76;  #10 
a = 8'd71; b = 8'd77;  #10 
a = 8'd71; b = 8'd78;  #10 
a = 8'd71; b = 8'd79;  #10 
a = 8'd71; b = 8'd80;  #10 
a = 8'd71; b = 8'd81;  #10 
a = 8'd71; b = 8'd82;  #10 
a = 8'd71; b = 8'd83;  #10 
a = 8'd71; b = 8'd84;  #10 
a = 8'd71; b = 8'd85;  #10 
a = 8'd71; b = 8'd86;  #10 
a = 8'd71; b = 8'd87;  #10 
a = 8'd71; b = 8'd88;  #10 
a = 8'd71; b = 8'd89;  #10 
a = 8'd71; b = 8'd90;  #10 
a = 8'd71; b = 8'd91;  #10 
a = 8'd71; b = 8'd92;  #10 
a = 8'd71; b = 8'd93;  #10 
a = 8'd71; b = 8'd94;  #10 
a = 8'd71; b = 8'd95;  #10 
a = 8'd71; b = 8'd96;  #10 
a = 8'd71; b = 8'd97;  #10 
a = 8'd71; b = 8'd98;  #10 
a = 8'd71; b = 8'd99;  #10 
a = 8'd71; b = 8'd100;  #10 
a = 8'd71; b = 8'd101;  #10 
a = 8'd71; b = 8'd102;  #10 
a = 8'd71; b = 8'd103;  #10 
a = 8'd71; b = 8'd104;  #10 
a = 8'd71; b = 8'd105;  #10 
a = 8'd71; b = 8'd106;  #10 
a = 8'd71; b = 8'd107;  #10 
a = 8'd71; b = 8'd108;  #10 
a = 8'd71; b = 8'd109;  #10 
a = 8'd71; b = 8'd110;  #10 
a = 8'd71; b = 8'd111;  #10 
a = 8'd71; b = 8'd112;  #10 
a = 8'd71; b = 8'd113;  #10 
a = 8'd71; b = 8'd114;  #10 
a = 8'd71; b = 8'd115;  #10 
a = 8'd71; b = 8'd116;  #10 
a = 8'd71; b = 8'd117;  #10 
a = 8'd71; b = 8'd118;  #10 
a = 8'd71; b = 8'd119;  #10 
a = 8'd71; b = 8'd120;  #10 
a = 8'd71; b = 8'd121;  #10 
a = 8'd71; b = 8'd122;  #10 
a = 8'd71; b = 8'd123;  #10 
a = 8'd71; b = 8'd124;  #10 
a = 8'd71; b = 8'd125;  #10 
a = 8'd71; b = 8'd126;  #10 
a = 8'd71; b = 8'd127;  #10 
a = 8'd71; b = 8'd128;  #10 
a = 8'd71; b = 8'd129;  #10 
a = 8'd71; b = 8'd130;  #10 
a = 8'd71; b = 8'd131;  #10 
a = 8'd71; b = 8'd132;  #10 
a = 8'd71; b = 8'd133;  #10 
a = 8'd71; b = 8'd134;  #10 
a = 8'd71; b = 8'd135;  #10 
a = 8'd71; b = 8'd136;  #10 
a = 8'd71; b = 8'd137;  #10 
a = 8'd71; b = 8'd138;  #10 
a = 8'd71; b = 8'd139;  #10 
a = 8'd71; b = 8'd140;  #10 
a = 8'd71; b = 8'd141;  #10 
a = 8'd71; b = 8'd142;  #10 
a = 8'd71; b = 8'd143;  #10 
a = 8'd71; b = 8'd144;  #10 
a = 8'd71; b = 8'd145;  #10 
a = 8'd71; b = 8'd146;  #10 
a = 8'd71; b = 8'd147;  #10 
a = 8'd71; b = 8'd148;  #10 
a = 8'd71; b = 8'd149;  #10 
a = 8'd71; b = 8'd150;  #10 
a = 8'd71; b = 8'd151;  #10 
a = 8'd71; b = 8'd152;  #10 
a = 8'd71; b = 8'd153;  #10 
a = 8'd71; b = 8'd154;  #10 
a = 8'd71; b = 8'd155;  #10 
a = 8'd71; b = 8'd156;  #10 
a = 8'd71; b = 8'd157;  #10 
a = 8'd71; b = 8'd158;  #10 
a = 8'd71; b = 8'd159;  #10 
a = 8'd71; b = 8'd160;  #10 
a = 8'd71; b = 8'd161;  #10 
a = 8'd71; b = 8'd162;  #10 
a = 8'd71; b = 8'd163;  #10 
a = 8'd71; b = 8'd164;  #10 
a = 8'd71; b = 8'd165;  #10 
a = 8'd71; b = 8'd166;  #10 
a = 8'd71; b = 8'd167;  #10 
a = 8'd71; b = 8'd168;  #10 
a = 8'd71; b = 8'd169;  #10 
a = 8'd71; b = 8'd170;  #10 
a = 8'd71; b = 8'd171;  #10 
a = 8'd71; b = 8'd172;  #10 
a = 8'd71; b = 8'd173;  #10 
a = 8'd71; b = 8'd174;  #10 
a = 8'd71; b = 8'd175;  #10 
a = 8'd71; b = 8'd176;  #10 
a = 8'd71; b = 8'd177;  #10 
a = 8'd71; b = 8'd178;  #10 
a = 8'd71; b = 8'd179;  #10 
a = 8'd71; b = 8'd180;  #10 
a = 8'd71; b = 8'd181;  #10 
a = 8'd71; b = 8'd182;  #10 
a = 8'd71; b = 8'd183;  #10 
a = 8'd71; b = 8'd184;  #10 
a = 8'd71; b = 8'd185;  #10 
a = 8'd71; b = 8'd186;  #10 
a = 8'd71; b = 8'd187;  #10 
a = 8'd71; b = 8'd188;  #10 
a = 8'd71; b = 8'd189;  #10 
a = 8'd71; b = 8'd190;  #10 
a = 8'd71; b = 8'd191;  #10 
a = 8'd71; b = 8'd192;  #10 
a = 8'd71; b = 8'd193;  #10 
a = 8'd71; b = 8'd194;  #10 
a = 8'd71; b = 8'd195;  #10 
a = 8'd71; b = 8'd196;  #10 
a = 8'd71; b = 8'd197;  #10 
a = 8'd71; b = 8'd198;  #10 
a = 8'd71; b = 8'd199;  #10 
a = 8'd71; b = 8'd200;  #10 
a = 8'd71; b = 8'd201;  #10 
a = 8'd71; b = 8'd202;  #10 
a = 8'd71; b = 8'd203;  #10 
a = 8'd71; b = 8'd204;  #10 
a = 8'd71; b = 8'd205;  #10 
a = 8'd71; b = 8'd206;  #10 
a = 8'd71; b = 8'd207;  #10 
a = 8'd71; b = 8'd208;  #10 
a = 8'd71; b = 8'd209;  #10 
a = 8'd71; b = 8'd210;  #10 
a = 8'd71; b = 8'd211;  #10 
a = 8'd71; b = 8'd212;  #10 
a = 8'd71; b = 8'd213;  #10 
a = 8'd71; b = 8'd214;  #10 
a = 8'd71; b = 8'd215;  #10 
a = 8'd71; b = 8'd216;  #10 
a = 8'd71; b = 8'd217;  #10 
a = 8'd71; b = 8'd218;  #10 
a = 8'd71; b = 8'd219;  #10 
a = 8'd71; b = 8'd220;  #10 
a = 8'd71; b = 8'd221;  #10 
a = 8'd71; b = 8'd222;  #10 
a = 8'd71; b = 8'd223;  #10 
a = 8'd71; b = 8'd224;  #10 
a = 8'd71; b = 8'd225;  #10 
a = 8'd71; b = 8'd226;  #10 
a = 8'd71; b = 8'd227;  #10 
a = 8'd71; b = 8'd228;  #10 
a = 8'd71; b = 8'd229;  #10 
a = 8'd71; b = 8'd230;  #10 
a = 8'd71; b = 8'd231;  #10 
a = 8'd71; b = 8'd232;  #10 
a = 8'd71; b = 8'd233;  #10 
a = 8'd71; b = 8'd234;  #10 
a = 8'd71; b = 8'd235;  #10 
a = 8'd71; b = 8'd236;  #10 
a = 8'd71; b = 8'd237;  #10 
a = 8'd71; b = 8'd238;  #10 
a = 8'd71; b = 8'd239;  #10 
a = 8'd71; b = 8'd240;  #10 
a = 8'd71; b = 8'd241;  #10 
a = 8'd71; b = 8'd242;  #10 
a = 8'd71; b = 8'd243;  #10 
a = 8'd71; b = 8'd244;  #10 
a = 8'd71; b = 8'd245;  #10 
a = 8'd71; b = 8'd246;  #10 
a = 8'd71; b = 8'd247;  #10 
a = 8'd71; b = 8'd248;  #10 
a = 8'd71; b = 8'd249;  #10 
a = 8'd71; b = 8'd250;  #10 
a = 8'd71; b = 8'd251;  #10 
a = 8'd71; b = 8'd252;  #10 
a = 8'd71; b = 8'd253;  #10 
a = 8'd71; b = 8'd254;  #10 
a = 8'd71; b = 8'd255;  #10 
a = 8'd72; b = 8'd0;  #10 
a = 8'd72; b = 8'd1;  #10 
a = 8'd72; b = 8'd2;  #10 
a = 8'd72; b = 8'd3;  #10 
a = 8'd72; b = 8'd4;  #10 
a = 8'd72; b = 8'd5;  #10 
a = 8'd72; b = 8'd6;  #10 
a = 8'd72; b = 8'd7;  #10 
a = 8'd72; b = 8'd8;  #10 
a = 8'd72; b = 8'd9;  #10 
a = 8'd72; b = 8'd10;  #10 
a = 8'd72; b = 8'd11;  #10 
a = 8'd72; b = 8'd12;  #10 
a = 8'd72; b = 8'd13;  #10 
a = 8'd72; b = 8'd14;  #10 
a = 8'd72; b = 8'd15;  #10 
a = 8'd72; b = 8'd16;  #10 
a = 8'd72; b = 8'd17;  #10 
a = 8'd72; b = 8'd18;  #10 
a = 8'd72; b = 8'd19;  #10 
a = 8'd72; b = 8'd20;  #10 
a = 8'd72; b = 8'd21;  #10 
a = 8'd72; b = 8'd22;  #10 
a = 8'd72; b = 8'd23;  #10 
a = 8'd72; b = 8'd24;  #10 
a = 8'd72; b = 8'd25;  #10 
a = 8'd72; b = 8'd26;  #10 
a = 8'd72; b = 8'd27;  #10 
a = 8'd72; b = 8'd28;  #10 
a = 8'd72; b = 8'd29;  #10 
a = 8'd72; b = 8'd30;  #10 
a = 8'd72; b = 8'd31;  #10 
a = 8'd72; b = 8'd32;  #10 
a = 8'd72; b = 8'd33;  #10 
a = 8'd72; b = 8'd34;  #10 
a = 8'd72; b = 8'd35;  #10 
a = 8'd72; b = 8'd36;  #10 
a = 8'd72; b = 8'd37;  #10 
a = 8'd72; b = 8'd38;  #10 
a = 8'd72; b = 8'd39;  #10 
a = 8'd72; b = 8'd40;  #10 
a = 8'd72; b = 8'd41;  #10 
a = 8'd72; b = 8'd42;  #10 
a = 8'd72; b = 8'd43;  #10 
a = 8'd72; b = 8'd44;  #10 
a = 8'd72; b = 8'd45;  #10 
a = 8'd72; b = 8'd46;  #10 
a = 8'd72; b = 8'd47;  #10 
a = 8'd72; b = 8'd48;  #10 
a = 8'd72; b = 8'd49;  #10 
a = 8'd72; b = 8'd50;  #10 
a = 8'd72; b = 8'd51;  #10 
a = 8'd72; b = 8'd52;  #10 
a = 8'd72; b = 8'd53;  #10 
a = 8'd72; b = 8'd54;  #10 
a = 8'd72; b = 8'd55;  #10 
a = 8'd72; b = 8'd56;  #10 
a = 8'd72; b = 8'd57;  #10 
a = 8'd72; b = 8'd58;  #10 
a = 8'd72; b = 8'd59;  #10 
a = 8'd72; b = 8'd60;  #10 
a = 8'd72; b = 8'd61;  #10 
a = 8'd72; b = 8'd62;  #10 
a = 8'd72; b = 8'd63;  #10 
a = 8'd72; b = 8'd64;  #10 
a = 8'd72; b = 8'd65;  #10 
a = 8'd72; b = 8'd66;  #10 
a = 8'd72; b = 8'd67;  #10 
a = 8'd72; b = 8'd68;  #10 
a = 8'd72; b = 8'd69;  #10 
a = 8'd72; b = 8'd70;  #10 
a = 8'd72; b = 8'd71;  #10 
a = 8'd72; b = 8'd72;  #10 
a = 8'd72; b = 8'd73;  #10 
a = 8'd72; b = 8'd74;  #10 
a = 8'd72; b = 8'd75;  #10 
a = 8'd72; b = 8'd76;  #10 
a = 8'd72; b = 8'd77;  #10 
a = 8'd72; b = 8'd78;  #10 
a = 8'd72; b = 8'd79;  #10 
a = 8'd72; b = 8'd80;  #10 
a = 8'd72; b = 8'd81;  #10 
a = 8'd72; b = 8'd82;  #10 
a = 8'd72; b = 8'd83;  #10 
a = 8'd72; b = 8'd84;  #10 
a = 8'd72; b = 8'd85;  #10 
a = 8'd72; b = 8'd86;  #10 
a = 8'd72; b = 8'd87;  #10 
a = 8'd72; b = 8'd88;  #10 
a = 8'd72; b = 8'd89;  #10 
a = 8'd72; b = 8'd90;  #10 
a = 8'd72; b = 8'd91;  #10 
a = 8'd72; b = 8'd92;  #10 
a = 8'd72; b = 8'd93;  #10 
a = 8'd72; b = 8'd94;  #10 
a = 8'd72; b = 8'd95;  #10 
a = 8'd72; b = 8'd96;  #10 
a = 8'd72; b = 8'd97;  #10 
a = 8'd72; b = 8'd98;  #10 
a = 8'd72; b = 8'd99;  #10 
a = 8'd72; b = 8'd100;  #10 
a = 8'd72; b = 8'd101;  #10 
a = 8'd72; b = 8'd102;  #10 
a = 8'd72; b = 8'd103;  #10 
a = 8'd72; b = 8'd104;  #10 
a = 8'd72; b = 8'd105;  #10 
a = 8'd72; b = 8'd106;  #10 
a = 8'd72; b = 8'd107;  #10 
a = 8'd72; b = 8'd108;  #10 
a = 8'd72; b = 8'd109;  #10 
a = 8'd72; b = 8'd110;  #10 
a = 8'd72; b = 8'd111;  #10 
a = 8'd72; b = 8'd112;  #10 
a = 8'd72; b = 8'd113;  #10 
a = 8'd72; b = 8'd114;  #10 
a = 8'd72; b = 8'd115;  #10 
a = 8'd72; b = 8'd116;  #10 
a = 8'd72; b = 8'd117;  #10 
a = 8'd72; b = 8'd118;  #10 
a = 8'd72; b = 8'd119;  #10 
a = 8'd72; b = 8'd120;  #10 
a = 8'd72; b = 8'd121;  #10 
a = 8'd72; b = 8'd122;  #10 
a = 8'd72; b = 8'd123;  #10 
a = 8'd72; b = 8'd124;  #10 
a = 8'd72; b = 8'd125;  #10 
a = 8'd72; b = 8'd126;  #10 
a = 8'd72; b = 8'd127;  #10 
a = 8'd72; b = 8'd128;  #10 
a = 8'd72; b = 8'd129;  #10 
a = 8'd72; b = 8'd130;  #10 
a = 8'd72; b = 8'd131;  #10 
a = 8'd72; b = 8'd132;  #10 
a = 8'd72; b = 8'd133;  #10 
a = 8'd72; b = 8'd134;  #10 
a = 8'd72; b = 8'd135;  #10 
a = 8'd72; b = 8'd136;  #10 
a = 8'd72; b = 8'd137;  #10 
a = 8'd72; b = 8'd138;  #10 
a = 8'd72; b = 8'd139;  #10 
a = 8'd72; b = 8'd140;  #10 
a = 8'd72; b = 8'd141;  #10 
a = 8'd72; b = 8'd142;  #10 
a = 8'd72; b = 8'd143;  #10 
a = 8'd72; b = 8'd144;  #10 
a = 8'd72; b = 8'd145;  #10 
a = 8'd72; b = 8'd146;  #10 
a = 8'd72; b = 8'd147;  #10 
a = 8'd72; b = 8'd148;  #10 
a = 8'd72; b = 8'd149;  #10 
a = 8'd72; b = 8'd150;  #10 
a = 8'd72; b = 8'd151;  #10 
a = 8'd72; b = 8'd152;  #10 
a = 8'd72; b = 8'd153;  #10 
a = 8'd72; b = 8'd154;  #10 
a = 8'd72; b = 8'd155;  #10 
a = 8'd72; b = 8'd156;  #10 
a = 8'd72; b = 8'd157;  #10 
a = 8'd72; b = 8'd158;  #10 
a = 8'd72; b = 8'd159;  #10 
a = 8'd72; b = 8'd160;  #10 
a = 8'd72; b = 8'd161;  #10 
a = 8'd72; b = 8'd162;  #10 
a = 8'd72; b = 8'd163;  #10 
a = 8'd72; b = 8'd164;  #10 
a = 8'd72; b = 8'd165;  #10 
a = 8'd72; b = 8'd166;  #10 
a = 8'd72; b = 8'd167;  #10 
a = 8'd72; b = 8'd168;  #10 
a = 8'd72; b = 8'd169;  #10 
a = 8'd72; b = 8'd170;  #10 
a = 8'd72; b = 8'd171;  #10 
a = 8'd72; b = 8'd172;  #10 
a = 8'd72; b = 8'd173;  #10 
a = 8'd72; b = 8'd174;  #10 
a = 8'd72; b = 8'd175;  #10 
a = 8'd72; b = 8'd176;  #10 
a = 8'd72; b = 8'd177;  #10 
a = 8'd72; b = 8'd178;  #10 
a = 8'd72; b = 8'd179;  #10 
a = 8'd72; b = 8'd180;  #10 
a = 8'd72; b = 8'd181;  #10 
a = 8'd72; b = 8'd182;  #10 
a = 8'd72; b = 8'd183;  #10 
a = 8'd72; b = 8'd184;  #10 
a = 8'd72; b = 8'd185;  #10 
a = 8'd72; b = 8'd186;  #10 
a = 8'd72; b = 8'd187;  #10 
a = 8'd72; b = 8'd188;  #10 
a = 8'd72; b = 8'd189;  #10 
a = 8'd72; b = 8'd190;  #10 
a = 8'd72; b = 8'd191;  #10 
a = 8'd72; b = 8'd192;  #10 
a = 8'd72; b = 8'd193;  #10 
a = 8'd72; b = 8'd194;  #10 
a = 8'd72; b = 8'd195;  #10 
a = 8'd72; b = 8'd196;  #10 
a = 8'd72; b = 8'd197;  #10 
a = 8'd72; b = 8'd198;  #10 
a = 8'd72; b = 8'd199;  #10 
a = 8'd72; b = 8'd200;  #10 
a = 8'd72; b = 8'd201;  #10 
a = 8'd72; b = 8'd202;  #10 
a = 8'd72; b = 8'd203;  #10 
a = 8'd72; b = 8'd204;  #10 
a = 8'd72; b = 8'd205;  #10 
a = 8'd72; b = 8'd206;  #10 
a = 8'd72; b = 8'd207;  #10 
a = 8'd72; b = 8'd208;  #10 
a = 8'd72; b = 8'd209;  #10 
a = 8'd72; b = 8'd210;  #10 
a = 8'd72; b = 8'd211;  #10 
a = 8'd72; b = 8'd212;  #10 
a = 8'd72; b = 8'd213;  #10 
a = 8'd72; b = 8'd214;  #10 
a = 8'd72; b = 8'd215;  #10 
a = 8'd72; b = 8'd216;  #10 
a = 8'd72; b = 8'd217;  #10 
a = 8'd72; b = 8'd218;  #10 
a = 8'd72; b = 8'd219;  #10 
a = 8'd72; b = 8'd220;  #10 
a = 8'd72; b = 8'd221;  #10 
a = 8'd72; b = 8'd222;  #10 
a = 8'd72; b = 8'd223;  #10 
a = 8'd72; b = 8'd224;  #10 
a = 8'd72; b = 8'd225;  #10 
a = 8'd72; b = 8'd226;  #10 
a = 8'd72; b = 8'd227;  #10 
a = 8'd72; b = 8'd228;  #10 
a = 8'd72; b = 8'd229;  #10 
a = 8'd72; b = 8'd230;  #10 
a = 8'd72; b = 8'd231;  #10 
a = 8'd72; b = 8'd232;  #10 
a = 8'd72; b = 8'd233;  #10 
a = 8'd72; b = 8'd234;  #10 
a = 8'd72; b = 8'd235;  #10 
a = 8'd72; b = 8'd236;  #10 
a = 8'd72; b = 8'd237;  #10 
a = 8'd72; b = 8'd238;  #10 
a = 8'd72; b = 8'd239;  #10 
a = 8'd72; b = 8'd240;  #10 
a = 8'd72; b = 8'd241;  #10 
a = 8'd72; b = 8'd242;  #10 
a = 8'd72; b = 8'd243;  #10 
a = 8'd72; b = 8'd244;  #10 
a = 8'd72; b = 8'd245;  #10 
a = 8'd72; b = 8'd246;  #10 
a = 8'd72; b = 8'd247;  #10 
a = 8'd72; b = 8'd248;  #10 
a = 8'd72; b = 8'd249;  #10 
a = 8'd72; b = 8'd250;  #10 
a = 8'd72; b = 8'd251;  #10 
a = 8'd72; b = 8'd252;  #10 
a = 8'd72; b = 8'd253;  #10 
a = 8'd72; b = 8'd254;  #10 
a = 8'd72; b = 8'd255;  #10 
a = 8'd73; b = 8'd0;  #10 
a = 8'd73; b = 8'd1;  #10 
a = 8'd73; b = 8'd2;  #10 
a = 8'd73; b = 8'd3;  #10 
a = 8'd73; b = 8'd4;  #10 
a = 8'd73; b = 8'd5;  #10 
a = 8'd73; b = 8'd6;  #10 
a = 8'd73; b = 8'd7;  #10 
a = 8'd73; b = 8'd8;  #10 
a = 8'd73; b = 8'd9;  #10 
a = 8'd73; b = 8'd10;  #10 
a = 8'd73; b = 8'd11;  #10 
a = 8'd73; b = 8'd12;  #10 
a = 8'd73; b = 8'd13;  #10 
a = 8'd73; b = 8'd14;  #10 
a = 8'd73; b = 8'd15;  #10 
a = 8'd73; b = 8'd16;  #10 
a = 8'd73; b = 8'd17;  #10 
a = 8'd73; b = 8'd18;  #10 
a = 8'd73; b = 8'd19;  #10 
a = 8'd73; b = 8'd20;  #10 
a = 8'd73; b = 8'd21;  #10 
a = 8'd73; b = 8'd22;  #10 
a = 8'd73; b = 8'd23;  #10 
a = 8'd73; b = 8'd24;  #10 
a = 8'd73; b = 8'd25;  #10 
a = 8'd73; b = 8'd26;  #10 
a = 8'd73; b = 8'd27;  #10 
a = 8'd73; b = 8'd28;  #10 
a = 8'd73; b = 8'd29;  #10 
a = 8'd73; b = 8'd30;  #10 
a = 8'd73; b = 8'd31;  #10 
a = 8'd73; b = 8'd32;  #10 
a = 8'd73; b = 8'd33;  #10 
a = 8'd73; b = 8'd34;  #10 
a = 8'd73; b = 8'd35;  #10 
a = 8'd73; b = 8'd36;  #10 
a = 8'd73; b = 8'd37;  #10 
a = 8'd73; b = 8'd38;  #10 
a = 8'd73; b = 8'd39;  #10 
a = 8'd73; b = 8'd40;  #10 
a = 8'd73; b = 8'd41;  #10 
a = 8'd73; b = 8'd42;  #10 
a = 8'd73; b = 8'd43;  #10 
a = 8'd73; b = 8'd44;  #10 
a = 8'd73; b = 8'd45;  #10 
a = 8'd73; b = 8'd46;  #10 
a = 8'd73; b = 8'd47;  #10 
a = 8'd73; b = 8'd48;  #10 
a = 8'd73; b = 8'd49;  #10 
a = 8'd73; b = 8'd50;  #10 
a = 8'd73; b = 8'd51;  #10 
a = 8'd73; b = 8'd52;  #10 
a = 8'd73; b = 8'd53;  #10 
a = 8'd73; b = 8'd54;  #10 
a = 8'd73; b = 8'd55;  #10 
a = 8'd73; b = 8'd56;  #10 
a = 8'd73; b = 8'd57;  #10 
a = 8'd73; b = 8'd58;  #10 
a = 8'd73; b = 8'd59;  #10 
a = 8'd73; b = 8'd60;  #10 
a = 8'd73; b = 8'd61;  #10 
a = 8'd73; b = 8'd62;  #10 
a = 8'd73; b = 8'd63;  #10 
a = 8'd73; b = 8'd64;  #10 
a = 8'd73; b = 8'd65;  #10 
a = 8'd73; b = 8'd66;  #10 
a = 8'd73; b = 8'd67;  #10 
a = 8'd73; b = 8'd68;  #10 
a = 8'd73; b = 8'd69;  #10 
a = 8'd73; b = 8'd70;  #10 
a = 8'd73; b = 8'd71;  #10 
a = 8'd73; b = 8'd72;  #10 
a = 8'd73; b = 8'd73;  #10 
a = 8'd73; b = 8'd74;  #10 
a = 8'd73; b = 8'd75;  #10 
a = 8'd73; b = 8'd76;  #10 
a = 8'd73; b = 8'd77;  #10 
a = 8'd73; b = 8'd78;  #10 
a = 8'd73; b = 8'd79;  #10 
a = 8'd73; b = 8'd80;  #10 
a = 8'd73; b = 8'd81;  #10 
a = 8'd73; b = 8'd82;  #10 
a = 8'd73; b = 8'd83;  #10 
a = 8'd73; b = 8'd84;  #10 
a = 8'd73; b = 8'd85;  #10 
a = 8'd73; b = 8'd86;  #10 
a = 8'd73; b = 8'd87;  #10 
a = 8'd73; b = 8'd88;  #10 
a = 8'd73; b = 8'd89;  #10 
a = 8'd73; b = 8'd90;  #10 
a = 8'd73; b = 8'd91;  #10 
a = 8'd73; b = 8'd92;  #10 
a = 8'd73; b = 8'd93;  #10 
a = 8'd73; b = 8'd94;  #10 
a = 8'd73; b = 8'd95;  #10 
a = 8'd73; b = 8'd96;  #10 
a = 8'd73; b = 8'd97;  #10 
a = 8'd73; b = 8'd98;  #10 
a = 8'd73; b = 8'd99;  #10 
a = 8'd73; b = 8'd100;  #10 
a = 8'd73; b = 8'd101;  #10 
a = 8'd73; b = 8'd102;  #10 
a = 8'd73; b = 8'd103;  #10 
a = 8'd73; b = 8'd104;  #10 
a = 8'd73; b = 8'd105;  #10 
a = 8'd73; b = 8'd106;  #10 
a = 8'd73; b = 8'd107;  #10 
a = 8'd73; b = 8'd108;  #10 
a = 8'd73; b = 8'd109;  #10 
a = 8'd73; b = 8'd110;  #10 
a = 8'd73; b = 8'd111;  #10 
a = 8'd73; b = 8'd112;  #10 
a = 8'd73; b = 8'd113;  #10 
a = 8'd73; b = 8'd114;  #10 
a = 8'd73; b = 8'd115;  #10 
a = 8'd73; b = 8'd116;  #10 
a = 8'd73; b = 8'd117;  #10 
a = 8'd73; b = 8'd118;  #10 
a = 8'd73; b = 8'd119;  #10 
a = 8'd73; b = 8'd120;  #10 
a = 8'd73; b = 8'd121;  #10 
a = 8'd73; b = 8'd122;  #10 
a = 8'd73; b = 8'd123;  #10 
a = 8'd73; b = 8'd124;  #10 
a = 8'd73; b = 8'd125;  #10 
a = 8'd73; b = 8'd126;  #10 
a = 8'd73; b = 8'd127;  #10 
a = 8'd73; b = 8'd128;  #10 
a = 8'd73; b = 8'd129;  #10 
a = 8'd73; b = 8'd130;  #10 
a = 8'd73; b = 8'd131;  #10 
a = 8'd73; b = 8'd132;  #10 
a = 8'd73; b = 8'd133;  #10 
a = 8'd73; b = 8'd134;  #10 
a = 8'd73; b = 8'd135;  #10 
a = 8'd73; b = 8'd136;  #10 
a = 8'd73; b = 8'd137;  #10 
a = 8'd73; b = 8'd138;  #10 
a = 8'd73; b = 8'd139;  #10 
a = 8'd73; b = 8'd140;  #10 
a = 8'd73; b = 8'd141;  #10 
a = 8'd73; b = 8'd142;  #10 
a = 8'd73; b = 8'd143;  #10 
a = 8'd73; b = 8'd144;  #10 
a = 8'd73; b = 8'd145;  #10 
a = 8'd73; b = 8'd146;  #10 
a = 8'd73; b = 8'd147;  #10 
a = 8'd73; b = 8'd148;  #10 
a = 8'd73; b = 8'd149;  #10 
a = 8'd73; b = 8'd150;  #10 
a = 8'd73; b = 8'd151;  #10 
a = 8'd73; b = 8'd152;  #10 
a = 8'd73; b = 8'd153;  #10 
a = 8'd73; b = 8'd154;  #10 
a = 8'd73; b = 8'd155;  #10 
a = 8'd73; b = 8'd156;  #10 
a = 8'd73; b = 8'd157;  #10 
a = 8'd73; b = 8'd158;  #10 
a = 8'd73; b = 8'd159;  #10 
a = 8'd73; b = 8'd160;  #10 
a = 8'd73; b = 8'd161;  #10 
a = 8'd73; b = 8'd162;  #10 
a = 8'd73; b = 8'd163;  #10 
a = 8'd73; b = 8'd164;  #10 
a = 8'd73; b = 8'd165;  #10 
a = 8'd73; b = 8'd166;  #10 
a = 8'd73; b = 8'd167;  #10 
a = 8'd73; b = 8'd168;  #10 
a = 8'd73; b = 8'd169;  #10 
a = 8'd73; b = 8'd170;  #10 
a = 8'd73; b = 8'd171;  #10 
a = 8'd73; b = 8'd172;  #10 
a = 8'd73; b = 8'd173;  #10 
a = 8'd73; b = 8'd174;  #10 
a = 8'd73; b = 8'd175;  #10 
a = 8'd73; b = 8'd176;  #10 
a = 8'd73; b = 8'd177;  #10 
a = 8'd73; b = 8'd178;  #10 
a = 8'd73; b = 8'd179;  #10 
a = 8'd73; b = 8'd180;  #10 
a = 8'd73; b = 8'd181;  #10 
a = 8'd73; b = 8'd182;  #10 
a = 8'd73; b = 8'd183;  #10 
a = 8'd73; b = 8'd184;  #10 
a = 8'd73; b = 8'd185;  #10 
a = 8'd73; b = 8'd186;  #10 
a = 8'd73; b = 8'd187;  #10 
a = 8'd73; b = 8'd188;  #10 
a = 8'd73; b = 8'd189;  #10 
a = 8'd73; b = 8'd190;  #10 
a = 8'd73; b = 8'd191;  #10 
a = 8'd73; b = 8'd192;  #10 
a = 8'd73; b = 8'd193;  #10 
a = 8'd73; b = 8'd194;  #10 
a = 8'd73; b = 8'd195;  #10 
a = 8'd73; b = 8'd196;  #10 
a = 8'd73; b = 8'd197;  #10 
a = 8'd73; b = 8'd198;  #10 
a = 8'd73; b = 8'd199;  #10 
a = 8'd73; b = 8'd200;  #10 
a = 8'd73; b = 8'd201;  #10 
a = 8'd73; b = 8'd202;  #10 
a = 8'd73; b = 8'd203;  #10 
a = 8'd73; b = 8'd204;  #10 
a = 8'd73; b = 8'd205;  #10 
a = 8'd73; b = 8'd206;  #10 
a = 8'd73; b = 8'd207;  #10 
a = 8'd73; b = 8'd208;  #10 
a = 8'd73; b = 8'd209;  #10 
a = 8'd73; b = 8'd210;  #10 
a = 8'd73; b = 8'd211;  #10 
a = 8'd73; b = 8'd212;  #10 
a = 8'd73; b = 8'd213;  #10 
a = 8'd73; b = 8'd214;  #10 
a = 8'd73; b = 8'd215;  #10 
a = 8'd73; b = 8'd216;  #10 
a = 8'd73; b = 8'd217;  #10 
a = 8'd73; b = 8'd218;  #10 
a = 8'd73; b = 8'd219;  #10 
a = 8'd73; b = 8'd220;  #10 
a = 8'd73; b = 8'd221;  #10 
a = 8'd73; b = 8'd222;  #10 
a = 8'd73; b = 8'd223;  #10 
a = 8'd73; b = 8'd224;  #10 
a = 8'd73; b = 8'd225;  #10 
a = 8'd73; b = 8'd226;  #10 
a = 8'd73; b = 8'd227;  #10 
a = 8'd73; b = 8'd228;  #10 
a = 8'd73; b = 8'd229;  #10 
a = 8'd73; b = 8'd230;  #10 
a = 8'd73; b = 8'd231;  #10 
a = 8'd73; b = 8'd232;  #10 
a = 8'd73; b = 8'd233;  #10 
a = 8'd73; b = 8'd234;  #10 
a = 8'd73; b = 8'd235;  #10 
a = 8'd73; b = 8'd236;  #10 
a = 8'd73; b = 8'd237;  #10 
a = 8'd73; b = 8'd238;  #10 
a = 8'd73; b = 8'd239;  #10 
a = 8'd73; b = 8'd240;  #10 
a = 8'd73; b = 8'd241;  #10 
a = 8'd73; b = 8'd242;  #10 
a = 8'd73; b = 8'd243;  #10 
a = 8'd73; b = 8'd244;  #10 
a = 8'd73; b = 8'd245;  #10 
a = 8'd73; b = 8'd246;  #10 
a = 8'd73; b = 8'd247;  #10 
a = 8'd73; b = 8'd248;  #10 
a = 8'd73; b = 8'd249;  #10 
a = 8'd73; b = 8'd250;  #10 
a = 8'd73; b = 8'd251;  #10 
a = 8'd73; b = 8'd252;  #10 
a = 8'd73; b = 8'd253;  #10 
a = 8'd73; b = 8'd254;  #10 
a = 8'd73; b = 8'd255;  #10 
a = 8'd74; b = 8'd0;  #10 
a = 8'd74; b = 8'd1;  #10 
a = 8'd74; b = 8'd2;  #10 
a = 8'd74; b = 8'd3;  #10 
a = 8'd74; b = 8'd4;  #10 
a = 8'd74; b = 8'd5;  #10 
a = 8'd74; b = 8'd6;  #10 
a = 8'd74; b = 8'd7;  #10 
a = 8'd74; b = 8'd8;  #10 
a = 8'd74; b = 8'd9;  #10 
a = 8'd74; b = 8'd10;  #10 
a = 8'd74; b = 8'd11;  #10 
a = 8'd74; b = 8'd12;  #10 
a = 8'd74; b = 8'd13;  #10 
a = 8'd74; b = 8'd14;  #10 
a = 8'd74; b = 8'd15;  #10 
a = 8'd74; b = 8'd16;  #10 
a = 8'd74; b = 8'd17;  #10 
a = 8'd74; b = 8'd18;  #10 
a = 8'd74; b = 8'd19;  #10 
a = 8'd74; b = 8'd20;  #10 
a = 8'd74; b = 8'd21;  #10 
a = 8'd74; b = 8'd22;  #10 
a = 8'd74; b = 8'd23;  #10 
a = 8'd74; b = 8'd24;  #10 
a = 8'd74; b = 8'd25;  #10 
a = 8'd74; b = 8'd26;  #10 
a = 8'd74; b = 8'd27;  #10 
a = 8'd74; b = 8'd28;  #10 
a = 8'd74; b = 8'd29;  #10 
a = 8'd74; b = 8'd30;  #10 
a = 8'd74; b = 8'd31;  #10 
a = 8'd74; b = 8'd32;  #10 
a = 8'd74; b = 8'd33;  #10 
a = 8'd74; b = 8'd34;  #10 
a = 8'd74; b = 8'd35;  #10 
a = 8'd74; b = 8'd36;  #10 
a = 8'd74; b = 8'd37;  #10 
a = 8'd74; b = 8'd38;  #10 
a = 8'd74; b = 8'd39;  #10 
a = 8'd74; b = 8'd40;  #10 
a = 8'd74; b = 8'd41;  #10 
a = 8'd74; b = 8'd42;  #10 
a = 8'd74; b = 8'd43;  #10 
a = 8'd74; b = 8'd44;  #10 
a = 8'd74; b = 8'd45;  #10 
a = 8'd74; b = 8'd46;  #10 
a = 8'd74; b = 8'd47;  #10 
a = 8'd74; b = 8'd48;  #10 
a = 8'd74; b = 8'd49;  #10 
a = 8'd74; b = 8'd50;  #10 
a = 8'd74; b = 8'd51;  #10 
a = 8'd74; b = 8'd52;  #10 
a = 8'd74; b = 8'd53;  #10 
a = 8'd74; b = 8'd54;  #10 
a = 8'd74; b = 8'd55;  #10 
a = 8'd74; b = 8'd56;  #10 
a = 8'd74; b = 8'd57;  #10 
a = 8'd74; b = 8'd58;  #10 
a = 8'd74; b = 8'd59;  #10 
a = 8'd74; b = 8'd60;  #10 
a = 8'd74; b = 8'd61;  #10 
a = 8'd74; b = 8'd62;  #10 
a = 8'd74; b = 8'd63;  #10 
a = 8'd74; b = 8'd64;  #10 
a = 8'd74; b = 8'd65;  #10 
a = 8'd74; b = 8'd66;  #10 
a = 8'd74; b = 8'd67;  #10 
a = 8'd74; b = 8'd68;  #10 
a = 8'd74; b = 8'd69;  #10 
a = 8'd74; b = 8'd70;  #10 
a = 8'd74; b = 8'd71;  #10 
a = 8'd74; b = 8'd72;  #10 
a = 8'd74; b = 8'd73;  #10 
a = 8'd74; b = 8'd74;  #10 
a = 8'd74; b = 8'd75;  #10 
a = 8'd74; b = 8'd76;  #10 
a = 8'd74; b = 8'd77;  #10 
a = 8'd74; b = 8'd78;  #10 
a = 8'd74; b = 8'd79;  #10 
a = 8'd74; b = 8'd80;  #10 
a = 8'd74; b = 8'd81;  #10 
a = 8'd74; b = 8'd82;  #10 
a = 8'd74; b = 8'd83;  #10 
a = 8'd74; b = 8'd84;  #10 
a = 8'd74; b = 8'd85;  #10 
a = 8'd74; b = 8'd86;  #10 
a = 8'd74; b = 8'd87;  #10 
a = 8'd74; b = 8'd88;  #10 
a = 8'd74; b = 8'd89;  #10 
a = 8'd74; b = 8'd90;  #10 
a = 8'd74; b = 8'd91;  #10 
a = 8'd74; b = 8'd92;  #10 
a = 8'd74; b = 8'd93;  #10 
a = 8'd74; b = 8'd94;  #10 
a = 8'd74; b = 8'd95;  #10 
a = 8'd74; b = 8'd96;  #10 
a = 8'd74; b = 8'd97;  #10 
a = 8'd74; b = 8'd98;  #10 
a = 8'd74; b = 8'd99;  #10 
a = 8'd74; b = 8'd100;  #10 
a = 8'd74; b = 8'd101;  #10 
a = 8'd74; b = 8'd102;  #10 
a = 8'd74; b = 8'd103;  #10 
a = 8'd74; b = 8'd104;  #10 
a = 8'd74; b = 8'd105;  #10 
a = 8'd74; b = 8'd106;  #10 
a = 8'd74; b = 8'd107;  #10 
a = 8'd74; b = 8'd108;  #10 
a = 8'd74; b = 8'd109;  #10 
a = 8'd74; b = 8'd110;  #10 
a = 8'd74; b = 8'd111;  #10 
a = 8'd74; b = 8'd112;  #10 
a = 8'd74; b = 8'd113;  #10 
a = 8'd74; b = 8'd114;  #10 
a = 8'd74; b = 8'd115;  #10 
a = 8'd74; b = 8'd116;  #10 
a = 8'd74; b = 8'd117;  #10 
a = 8'd74; b = 8'd118;  #10 
a = 8'd74; b = 8'd119;  #10 
a = 8'd74; b = 8'd120;  #10 
a = 8'd74; b = 8'd121;  #10 
a = 8'd74; b = 8'd122;  #10 
a = 8'd74; b = 8'd123;  #10 
a = 8'd74; b = 8'd124;  #10 
a = 8'd74; b = 8'd125;  #10 
a = 8'd74; b = 8'd126;  #10 
a = 8'd74; b = 8'd127;  #10 
a = 8'd74; b = 8'd128;  #10 
a = 8'd74; b = 8'd129;  #10 
a = 8'd74; b = 8'd130;  #10 
a = 8'd74; b = 8'd131;  #10 
a = 8'd74; b = 8'd132;  #10 
a = 8'd74; b = 8'd133;  #10 
a = 8'd74; b = 8'd134;  #10 
a = 8'd74; b = 8'd135;  #10 
a = 8'd74; b = 8'd136;  #10 
a = 8'd74; b = 8'd137;  #10 
a = 8'd74; b = 8'd138;  #10 
a = 8'd74; b = 8'd139;  #10 
a = 8'd74; b = 8'd140;  #10 
a = 8'd74; b = 8'd141;  #10 
a = 8'd74; b = 8'd142;  #10 
a = 8'd74; b = 8'd143;  #10 
a = 8'd74; b = 8'd144;  #10 
a = 8'd74; b = 8'd145;  #10 
a = 8'd74; b = 8'd146;  #10 
a = 8'd74; b = 8'd147;  #10 
a = 8'd74; b = 8'd148;  #10 
a = 8'd74; b = 8'd149;  #10 
a = 8'd74; b = 8'd150;  #10 
a = 8'd74; b = 8'd151;  #10 
a = 8'd74; b = 8'd152;  #10 
a = 8'd74; b = 8'd153;  #10 
a = 8'd74; b = 8'd154;  #10 
a = 8'd74; b = 8'd155;  #10 
a = 8'd74; b = 8'd156;  #10 
a = 8'd74; b = 8'd157;  #10 
a = 8'd74; b = 8'd158;  #10 
a = 8'd74; b = 8'd159;  #10 
a = 8'd74; b = 8'd160;  #10 
a = 8'd74; b = 8'd161;  #10 
a = 8'd74; b = 8'd162;  #10 
a = 8'd74; b = 8'd163;  #10 
a = 8'd74; b = 8'd164;  #10 
a = 8'd74; b = 8'd165;  #10 
a = 8'd74; b = 8'd166;  #10 
a = 8'd74; b = 8'd167;  #10 
a = 8'd74; b = 8'd168;  #10 
a = 8'd74; b = 8'd169;  #10 
a = 8'd74; b = 8'd170;  #10 
a = 8'd74; b = 8'd171;  #10 
a = 8'd74; b = 8'd172;  #10 
a = 8'd74; b = 8'd173;  #10 
a = 8'd74; b = 8'd174;  #10 
a = 8'd74; b = 8'd175;  #10 
a = 8'd74; b = 8'd176;  #10 
a = 8'd74; b = 8'd177;  #10 
a = 8'd74; b = 8'd178;  #10 
a = 8'd74; b = 8'd179;  #10 
a = 8'd74; b = 8'd180;  #10 
a = 8'd74; b = 8'd181;  #10 
a = 8'd74; b = 8'd182;  #10 
a = 8'd74; b = 8'd183;  #10 
a = 8'd74; b = 8'd184;  #10 
a = 8'd74; b = 8'd185;  #10 
a = 8'd74; b = 8'd186;  #10 
a = 8'd74; b = 8'd187;  #10 
a = 8'd74; b = 8'd188;  #10 
a = 8'd74; b = 8'd189;  #10 
a = 8'd74; b = 8'd190;  #10 
a = 8'd74; b = 8'd191;  #10 
a = 8'd74; b = 8'd192;  #10 
a = 8'd74; b = 8'd193;  #10 
a = 8'd74; b = 8'd194;  #10 
a = 8'd74; b = 8'd195;  #10 
a = 8'd74; b = 8'd196;  #10 
a = 8'd74; b = 8'd197;  #10 
a = 8'd74; b = 8'd198;  #10 
a = 8'd74; b = 8'd199;  #10 
a = 8'd74; b = 8'd200;  #10 
a = 8'd74; b = 8'd201;  #10 
a = 8'd74; b = 8'd202;  #10 
a = 8'd74; b = 8'd203;  #10 
a = 8'd74; b = 8'd204;  #10 
a = 8'd74; b = 8'd205;  #10 
a = 8'd74; b = 8'd206;  #10 
a = 8'd74; b = 8'd207;  #10 
a = 8'd74; b = 8'd208;  #10 
a = 8'd74; b = 8'd209;  #10 
a = 8'd74; b = 8'd210;  #10 
a = 8'd74; b = 8'd211;  #10 
a = 8'd74; b = 8'd212;  #10 
a = 8'd74; b = 8'd213;  #10 
a = 8'd74; b = 8'd214;  #10 
a = 8'd74; b = 8'd215;  #10 
a = 8'd74; b = 8'd216;  #10 
a = 8'd74; b = 8'd217;  #10 
a = 8'd74; b = 8'd218;  #10 
a = 8'd74; b = 8'd219;  #10 
a = 8'd74; b = 8'd220;  #10 
a = 8'd74; b = 8'd221;  #10 
a = 8'd74; b = 8'd222;  #10 
a = 8'd74; b = 8'd223;  #10 
a = 8'd74; b = 8'd224;  #10 
a = 8'd74; b = 8'd225;  #10 
a = 8'd74; b = 8'd226;  #10 
a = 8'd74; b = 8'd227;  #10 
a = 8'd74; b = 8'd228;  #10 
a = 8'd74; b = 8'd229;  #10 
a = 8'd74; b = 8'd230;  #10 
a = 8'd74; b = 8'd231;  #10 
a = 8'd74; b = 8'd232;  #10 
a = 8'd74; b = 8'd233;  #10 
a = 8'd74; b = 8'd234;  #10 
a = 8'd74; b = 8'd235;  #10 
a = 8'd74; b = 8'd236;  #10 
a = 8'd74; b = 8'd237;  #10 
a = 8'd74; b = 8'd238;  #10 
a = 8'd74; b = 8'd239;  #10 
a = 8'd74; b = 8'd240;  #10 
a = 8'd74; b = 8'd241;  #10 
a = 8'd74; b = 8'd242;  #10 
a = 8'd74; b = 8'd243;  #10 
a = 8'd74; b = 8'd244;  #10 
a = 8'd74; b = 8'd245;  #10 
a = 8'd74; b = 8'd246;  #10 
a = 8'd74; b = 8'd247;  #10 
a = 8'd74; b = 8'd248;  #10 
a = 8'd74; b = 8'd249;  #10 
a = 8'd74; b = 8'd250;  #10 
a = 8'd74; b = 8'd251;  #10 
a = 8'd74; b = 8'd252;  #10 
a = 8'd74; b = 8'd253;  #10 
a = 8'd74; b = 8'd254;  #10 
a = 8'd74; b = 8'd255;  #10 
a = 8'd75; b = 8'd0;  #10 
a = 8'd75; b = 8'd1;  #10 
a = 8'd75; b = 8'd2;  #10 
a = 8'd75; b = 8'd3;  #10 
a = 8'd75; b = 8'd4;  #10 
a = 8'd75; b = 8'd5;  #10 
a = 8'd75; b = 8'd6;  #10 
a = 8'd75; b = 8'd7;  #10 
a = 8'd75; b = 8'd8;  #10 
a = 8'd75; b = 8'd9;  #10 
a = 8'd75; b = 8'd10;  #10 
a = 8'd75; b = 8'd11;  #10 
a = 8'd75; b = 8'd12;  #10 
a = 8'd75; b = 8'd13;  #10 
a = 8'd75; b = 8'd14;  #10 
a = 8'd75; b = 8'd15;  #10 
a = 8'd75; b = 8'd16;  #10 
a = 8'd75; b = 8'd17;  #10 
a = 8'd75; b = 8'd18;  #10 
a = 8'd75; b = 8'd19;  #10 
a = 8'd75; b = 8'd20;  #10 
a = 8'd75; b = 8'd21;  #10 
a = 8'd75; b = 8'd22;  #10 
a = 8'd75; b = 8'd23;  #10 
a = 8'd75; b = 8'd24;  #10 
a = 8'd75; b = 8'd25;  #10 
a = 8'd75; b = 8'd26;  #10 
a = 8'd75; b = 8'd27;  #10 
a = 8'd75; b = 8'd28;  #10 
a = 8'd75; b = 8'd29;  #10 
a = 8'd75; b = 8'd30;  #10 
a = 8'd75; b = 8'd31;  #10 
a = 8'd75; b = 8'd32;  #10 
a = 8'd75; b = 8'd33;  #10 
a = 8'd75; b = 8'd34;  #10 
a = 8'd75; b = 8'd35;  #10 
a = 8'd75; b = 8'd36;  #10 
a = 8'd75; b = 8'd37;  #10 
a = 8'd75; b = 8'd38;  #10 
a = 8'd75; b = 8'd39;  #10 
a = 8'd75; b = 8'd40;  #10 
a = 8'd75; b = 8'd41;  #10 
a = 8'd75; b = 8'd42;  #10 
a = 8'd75; b = 8'd43;  #10 
a = 8'd75; b = 8'd44;  #10 
a = 8'd75; b = 8'd45;  #10 
a = 8'd75; b = 8'd46;  #10 
a = 8'd75; b = 8'd47;  #10 
a = 8'd75; b = 8'd48;  #10 
a = 8'd75; b = 8'd49;  #10 
a = 8'd75; b = 8'd50;  #10 
a = 8'd75; b = 8'd51;  #10 
a = 8'd75; b = 8'd52;  #10 
a = 8'd75; b = 8'd53;  #10 
a = 8'd75; b = 8'd54;  #10 
a = 8'd75; b = 8'd55;  #10 
a = 8'd75; b = 8'd56;  #10 
a = 8'd75; b = 8'd57;  #10 
a = 8'd75; b = 8'd58;  #10 
a = 8'd75; b = 8'd59;  #10 
a = 8'd75; b = 8'd60;  #10 
a = 8'd75; b = 8'd61;  #10 
a = 8'd75; b = 8'd62;  #10 
a = 8'd75; b = 8'd63;  #10 
a = 8'd75; b = 8'd64;  #10 
a = 8'd75; b = 8'd65;  #10 
a = 8'd75; b = 8'd66;  #10 
a = 8'd75; b = 8'd67;  #10 
a = 8'd75; b = 8'd68;  #10 
a = 8'd75; b = 8'd69;  #10 
a = 8'd75; b = 8'd70;  #10 
a = 8'd75; b = 8'd71;  #10 
a = 8'd75; b = 8'd72;  #10 
a = 8'd75; b = 8'd73;  #10 
a = 8'd75; b = 8'd74;  #10 
a = 8'd75; b = 8'd75;  #10 
a = 8'd75; b = 8'd76;  #10 
a = 8'd75; b = 8'd77;  #10 
a = 8'd75; b = 8'd78;  #10 
a = 8'd75; b = 8'd79;  #10 
a = 8'd75; b = 8'd80;  #10 
a = 8'd75; b = 8'd81;  #10 
a = 8'd75; b = 8'd82;  #10 
a = 8'd75; b = 8'd83;  #10 
a = 8'd75; b = 8'd84;  #10 
a = 8'd75; b = 8'd85;  #10 
a = 8'd75; b = 8'd86;  #10 
a = 8'd75; b = 8'd87;  #10 
a = 8'd75; b = 8'd88;  #10 
a = 8'd75; b = 8'd89;  #10 
a = 8'd75; b = 8'd90;  #10 
a = 8'd75; b = 8'd91;  #10 
a = 8'd75; b = 8'd92;  #10 
a = 8'd75; b = 8'd93;  #10 
a = 8'd75; b = 8'd94;  #10 
a = 8'd75; b = 8'd95;  #10 
a = 8'd75; b = 8'd96;  #10 
a = 8'd75; b = 8'd97;  #10 
a = 8'd75; b = 8'd98;  #10 
a = 8'd75; b = 8'd99;  #10 
a = 8'd75; b = 8'd100;  #10 
a = 8'd75; b = 8'd101;  #10 
a = 8'd75; b = 8'd102;  #10 
a = 8'd75; b = 8'd103;  #10 
a = 8'd75; b = 8'd104;  #10 
a = 8'd75; b = 8'd105;  #10 
a = 8'd75; b = 8'd106;  #10 
a = 8'd75; b = 8'd107;  #10 
a = 8'd75; b = 8'd108;  #10 
a = 8'd75; b = 8'd109;  #10 
a = 8'd75; b = 8'd110;  #10 
a = 8'd75; b = 8'd111;  #10 
a = 8'd75; b = 8'd112;  #10 
a = 8'd75; b = 8'd113;  #10 
a = 8'd75; b = 8'd114;  #10 
a = 8'd75; b = 8'd115;  #10 
a = 8'd75; b = 8'd116;  #10 
a = 8'd75; b = 8'd117;  #10 
a = 8'd75; b = 8'd118;  #10 
a = 8'd75; b = 8'd119;  #10 
a = 8'd75; b = 8'd120;  #10 
a = 8'd75; b = 8'd121;  #10 
a = 8'd75; b = 8'd122;  #10 
a = 8'd75; b = 8'd123;  #10 
a = 8'd75; b = 8'd124;  #10 
a = 8'd75; b = 8'd125;  #10 
a = 8'd75; b = 8'd126;  #10 
a = 8'd75; b = 8'd127;  #10 
a = 8'd75; b = 8'd128;  #10 
a = 8'd75; b = 8'd129;  #10 
a = 8'd75; b = 8'd130;  #10 
a = 8'd75; b = 8'd131;  #10 
a = 8'd75; b = 8'd132;  #10 
a = 8'd75; b = 8'd133;  #10 
a = 8'd75; b = 8'd134;  #10 
a = 8'd75; b = 8'd135;  #10 
a = 8'd75; b = 8'd136;  #10 
a = 8'd75; b = 8'd137;  #10 
a = 8'd75; b = 8'd138;  #10 
a = 8'd75; b = 8'd139;  #10 
a = 8'd75; b = 8'd140;  #10 
a = 8'd75; b = 8'd141;  #10 
a = 8'd75; b = 8'd142;  #10 
a = 8'd75; b = 8'd143;  #10 
a = 8'd75; b = 8'd144;  #10 
a = 8'd75; b = 8'd145;  #10 
a = 8'd75; b = 8'd146;  #10 
a = 8'd75; b = 8'd147;  #10 
a = 8'd75; b = 8'd148;  #10 
a = 8'd75; b = 8'd149;  #10 
a = 8'd75; b = 8'd150;  #10 
a = 8'd75; b = 8'd151;  #10 
a = 8'd75; b = 8'd152;  #10 
a = 8'd75; b = 8'd153;  #10 
a = 8'd75; b = 8'd154;  #10 
a = 8'd75; b = 8'd155;  #10 
a = 8'd75; b = 8'd156;  #10 
a = 8'd75; b = 8'd157;  #10 
a = 8'd75; b = 8'd158;  #10 
a = 8'd75; b = 8'd159;  #10 
a = 8'd75; b = 8'd160;  #10 
a = 8'd75; b = 8'd161;  #10 
a = 8'd75; b = 8'd162;  #10 
a = 8'd75; b = 8'd163;  #10 
a = 8'd75; b = 8'd164;  #10 
a = 8'd75; b = 8'd165;  #10 
a = 8'd75; b = 8'd166;  #10 
a = 8'd75; b = 8'd167;  #10 
a = 8'd75; b = 8'd168;  #10 
a = 8'd75; b = 8'd169;  #10 
a = 8'd75; b = 8'd170;  #10 
a = 8'd75; b = 8'd171;  #10 
a = 8'd75; b = 8'd172;  #10 
a = 8'd75; b = 8'd173;  #10 
a = 8'd75; b = 8'd174;  #10 
a = 8'd75; b = 8'd175;  #10 
a = 8'd75; b = 8'd176;  #10 
a = 8'd75; b = 8'd177;  #10 
a = 8'd75; b = 8'd178;  #10 
a = 8'd75; b = 8'd179;  #10 
a = 8'd75; b = 8'd180;  #10 
a = 8'd75; b = 8'd181;  #10 
a = 8'd75; b = 8'd182;  #10 
a = 8'd75; b = 8'd183;  #10 
a = 8'd75; b = 8'd184;  #10 
a = 8'd75; b = 8'd185;  #10 
a = 8'd75; b = 8'd186;  #10 
a = 8'd75; b = 8'd187;  #10 
a = 8'd75; b = 8'd188;  #10 
a = 8'd75; b = 8'd189;  #10 
a = 8'd75; b = 8'd190;  #10 
a = 8'd75; b = 8'd191;  #10 
a = 8'd75; b = 8'd192;  #10 
a = 8'd75; b = 8'd193;  #10 
a = 8'd75; b = 8'd194;  #10 
a = 8'd75; b = 8'd195;  #10 
a = 8'd75; b = 8'd196;  #10 
a = 8'd75; b = 8'd197;  #10 
a = 8'd75; b = 8'd198;  #10 
a = 8'd75; b = 8'd199;  #10 
a = 8'd75; b = 8'd200;  #10 
a = 8'd75; b = 8'd201;  #10 
a = 8'd75; b = 8'd202;  #10 
a = 8'd75; b = 8'd203;  #10 
a = 8'd75; b = 8'd204;  #10 
a = 8'd75; b = 8'd205;  #10 
a = 8'd75; b = 8'd206;  #10 
a = 8'd75; b = 8'd207;  #10 
a = 8'd75; b = 8'd208;  #10 
a = 8'd75; b = 8'd209;  #10 
a = 8'd75; b = 8'd210;  #10 
a = 8'd75; b = 8'd211;  #10 
a = 8'd75; b = 8'd212;  #10 
a = 8'd75; b = 8'd213;  #10 
a = 8'd75; b = 8'd214;  #10 
a = 8'd75; b = 8'd215;  #10 
a = 8'd75; b = 8'd216;  #10 
a = 8'd75; b = 8'd217;  #10 
a = 8'd75; b = 8'd218;  #10 
a = 8'd75; b = 8'd219;  #10 
a = 8'd75; b = 8'd220;  #10 
a = 8'd75; b = 8'd221;  #10 
a = 8'd75; b = 8'd222;  #10 
a = 8'd75; b = 8'd223;  #10 
a = 8'd75; b = 8'd224;  #10 
a = 8'd75; b = 8'd225;  #10 
a = 8'd75; b = 8'd226;  #10 
a = 8'd75; b = 8'd227;  #10 
a = 8'd75; b = 8'd228;  #10 
a = 8'd75; b = 8'd229;  #10 
a = 8'd75; b = 8'd230;  #10 
a = 8'd75; b = 8'd231;  #10 
a = 8'd75; b = 8'd232;  #10 
a = 8'd75; b = 8'd233;  #10 
a = 8'd75; b = 8'd234;  #10 
a = 8'd75; b = 8'd235;  #10 
a = 8'd75; b = 8'd236;  #10 
a = 8'd75; b = 8'd237;  #10 
a = 8'd75; b = 8'd238;  #10 
a = 8'd75; b = 8'd239;  #10 
a = 8'd75; b = 8'd240;  #10 
a = 8'd75; b = 8'd241;  #10 
a = 8'd75; b = 8'd242;  #10 
a = 8'd75; b = 8'd243;  #10 
a = 8'd75; b = 8'd244;  #10 
a = 8'd75; b = 8'd245;  #10 
a = 8'd75; b = 8'd246;  #10 
a = 8'd75; b = 8'd247;  #10 
a = 8'd75; b = 8'd248;  #10 
a = 8'd75; b = 8'd249;  #10 
a = 8'd75; b = 8'd250;  #10 
a = 8'd75; b = 8'd251;  #10 
a = 8'd75; b = 8'd252;  #10 
a = 8'd75; b = 8'd253;  #10 
a = 8'd75; b = 8'd254;  #10 
a = 8'd75; b = 8'd255;  #10 
a = 8'd76; b = 8'd0;  #10 
a = 8'd76; b = 8'd1;  #10 
a = 8'd76; b = 8'd2;  #10 
a = 8'd76; b = 8'd3;  #10 
a = 8'd76; b = 8'd4;  #10 
a = 8'd76; b = 8'd5;  #10 
a = 8'd76; b = 8'd6;  #10 
a = 8'd76; b = 8'd7;  #10 
a = 8'd76; b = 8'd8;  #10 
a = 8'd76; b = 8'd9;  #10 
a = 8'd76; b = 8'd10;  #10 
a = 8'd76; b = 8'd11;  #10 
a = 8'd76; b = 8'd12;  #10 
a = 8'd76; b = 8'd13;  #10 
a = 8'd76; b = 8'd14;  #10 
a = 8'd76; b = 8'd15;  #10 
a = 8'd76; b = 8'd16;  #10 
a = 8'd76; b = 8'd17;  #10 
a = 8'd76; b = 8'd18;  #10 
a = 8'd76; b = 8'd19;  #10 
a = 8'd76; b = 8'd20;  #10 
a = 8'd76; b = 8'd21;  #10 
a = 8'd76; b = 8'd22;  #10 
a = 8'd76; b = 8'd23;  #10 
a = 8'd76; b = 8'd24;  #10 
a = 8'd76; b = 8'd25;  #10 
a = 8'd76; b = 8'd26;  #10 
a = 8'd76; b = 8'd27;  #10 
a = 8'd76; b = 8'd28;  #10 
a = 8'd76; b = 8'd29;  #10 
a = 8'd76; b = 8'd30;  #10 
a = 8'd76; b = 8'd31;  #10 
a = 8'd76; b = 8'd32;  #10 
a = 8'd76; b = 8'd33;  #10 
a = 8'd76; b = 8'd34;  #10 
a = 8'd76; b = 8'd35;  #10 
a = 8'd76; b = 8'd36;  #10 
a = 8'd76; b = 8'd37;  #10 
a = 8'd76; b = 8'd38;  #10 
a = 8'd76; b = 8'd39;  #10 
a = 8'd76; b = 8'd40;  #10 
a = 8'd76; b = 8'd41;  #10 
a = 8'd76; b = 8'd42;  #10 
a = 8'd76; b = 8'd43;  #10 
a = 8'd76; b = 8'd44;  #10 
a = 8'd76; b = 8'd45;  #10 
a = 8'd76; b = 8'd46;  #10 
a = 8'd76; b = 8'd47;  #10 
a = 8'd76; b = 8'd48;  #10 
a = 8'd76; b = 8'd49;  #10 
a = 8'd76; b = 8'd50;  #10 
a = 8'd76; b = 8'd51;  #10 
a = 8'd76; b = 8'd52;  #10 
a = 8'd76; b = 8'd53;  #10 
a = 8'd76; b = 8'd54;  #10 
a = 8'd76; b = 8'd55;  #10 
a = 8'd76; b = 8'd56;  #10 
a = 8'd76; b = 8'd57;  #10 
a = 8'd76; b = 8'd58;  #10 
a = 8'd76; b = 8'd59;  #10 
a = 8'd76; b = 8'd60;  #10 
a = 8'd76; b = 8'd61;  #10 
a = 8'd76; b = 8'd62;  #10 
a = 8'd76; b = 8'd63;  #10 
a = 8'd76; b = 8'd64;  #10 
a = 8'd76; b = 8'd65;  #10 
a = 8'd76; b = 8'd66;  #10 
a = 8'd76; b = 8'd67;  #10 
a = 8'd76; b = 8'd68;  #10 
a = 8'd76; b = 8'd69;  #10 
a = 8'd76; b = 8'd70;  #10 
a = 8'd76; b = 8'd71;  #10 
a = 8'd76; b = 8'd72;  #10 
a = 8'd76; b = 8'd73;  #10 
a = 8'd76; b = 8'd74;  #10 
a = 8'd76; b = 8'd75;  #10 
a = 8'd76; b = 8'd76;  #10 
a = 8'd76; b = 8'd77;  #10 
a = 8'd76; b = 8'd78;  #10 
a = 8'd76; b = 8'd79;  #10 
a = 8'd76; b = 8'd80;  #10 
a = 8'd76; b = 8'd81;  #10 
a = 8'd76; b = 8'd82;  #10 
a = 8'd76; b = 8'd83;  #10 
a = 8'd76; b = 8'd84;  #10 
a = 8'd76; b = 8'd85;  #10 
a = 8'd76; b = 8'd86;  #10 
a = 8'd76; b = 8'd87;  #10 
a = 8'd76; b = 8'd88;  #10 
a = 8'd76; b = 8'd89;  #10 
a = 8'd76; b = 8'd90;  #10 
a = 8'd76; b = 8'd91;  #10 
a = 8'd76; b = 8'd92;  #10 
a = 8'd76; b = 8'd93;  #10 
a = 8'd76; b = 8'd94;  #10 
a = 8'd76; b = 8'd95;  #10 
a = 8'd76; b = 8'd96;  #10 
a = 8'd76; b = 8'd97;  #10 
a = 8'd76; b = 8'd98;  #10 
a = 8'd76; b = 8'd99;  #10 
a = 8'd76; b = 8'd100;  #10 
a = 8'd76; b = 8'd101;  #10 
a = 8'd76; b = 8'd102;  #10 
a = 8'd76; b = 8'd103;  #10 
a = 8'd76; b = 8'd104;  #10 
a = 8'd76; b = 8'd105;  #10 
a = 8'd76; b = 8'd106;  #10 
a = 8'd76; b = 8'd107;  #10 
a = 8'd76; b = 8'd108;  #10 
a = 8'd76; b = 8'd109;  #10 
a = 8'd76; b = 8'd110;  #10 
a = 8'd76; b = 8'd111;  #10 
a = 8'd76; b = 8'd112;  #10 
a = 8'd76; b = 8'd113;  #10 
a = 8'd76; b = 8'd114;  #10 
a = 8'd76; b = 8'd115;  #10 
a = 8'd76; b = 8'd116;  #10 
a = 8'd76; b = 8'd117;  #10 
a = 8'd76; b = 8'd118;  #10 
a = 8'd76; b = 8'd119;  #10 
a = 8'd76; b = 8'd120;  #10 
a = 8'd76; b = 8'd121;  #10 
a = 8'd76; b = 8'd122;  #10 
a = 8'd76; b = 8'd123;  #10 
a = 8'd76; b = 8'd124;  #10 
a = 8'd76; b = 8'd125;  #10 
a = 8'd76; b = 8'd126;  #10 
a = 8'd76; b = 8'd127;  #10 
a = 8'd76; b = 8'd128;  #10 
a = 8'd76; b = 8'd129;  #10 
a = 8'd76; b = 8'd130;  #10 
a = 8'd76; b = 8'd131;  #10 
a = 8'd76; b = 8'd132;  #10 
a = 8'd76; b = 8'd133;  #10 
a = 8'd76; b = 8'd134;  #10 
a = 8'd76; b = 8'd135;  #10 
a = 8'd76; b = 8'd136;  #10 
a = 8'd76; b = 8'd137;  #10 
a = 8'd76; b = 8'd138;  #10 
a = 8'd76; b = 8'd139;  #10 
a = 8'd76; b = 8'd140;  #10 
a = 8'd76; b = 8'd141;  #10 
a = 8'd76; b = 8'd142;  #10 
a = 8'd76; b = 8'd143;  #10 
a = 8'd76; b = 8'd144;  #10 
a = 8'd76; b = 8'd145;  #10 
a = 8'd76; b = 8'd146;  #10 
a = 8'd76; b = 8'd147;  #10 
a = 8'd76; b = 8'd148;  #10 
a = 8'd76; b = 8'd149;  #10 
a = 8'd76; b = 8'd150;  #10 
a = 8'd76; b = 8'd151;  #10 
a = 8'd76; b = 8'd152;  #10 
a = 8'd76; b = 8'd153;  #10 
a = 8'd76; b = 8'd154;  #10 
a = 8'd76; b = 8'd155;  #10 
a = 8'd76; b = 8'd156;  #10 
a = 8'd76; b = 8'd157;  #10 
a = 8'd76; b = 8'd158;  #10 
a = 8'd76; b = 8'd159;  #10 
a = 8'd76; b = 8'd160;  #10 
a = 8'd76; b = 8'd161;  #10 
a = 8'd76; b = 8'd162;  #10 
a = 8'd76; b = 8'd163;  #10 
a = 8'd76; b = 8'd164;  #10 
a = 8'd76; b = 8'd165;  #10 
a = 8'd76; b = 8'd166;  #10 
a = 8'd76; b = 8'd167;  #10 
a = 8'd76; b = 8'd168;  #10 
a = 8'd76; b = 8'd169;  #10 
a = 8'd76; b = 8'd170;  #10 
a = 8'd76; b = 8'd171;  #10 
a = 8'd76; b = 8'd172;  #10 
a = 8'd76; b = 8'd173;  #10 
a = 8'd76; b = 8'd174;  #10 
a = 8'd76; b = 8'd175;  #10 
a = 8'd76; b = 8'd176;  #10 
a = 8'd76; b = 8'd177;  #10 
a = 8'd76; b = 8'd178;  #10 
a = 8'd76; b = 8'd179;  #10 
a = 8'd76; b = 8'd180;  #10 
a = 8'd76; b = 8'd181;  #10 
a = 8'd76; b = 8'd182;  #10 
a = 8'd76; b = 8'd183;  #10 
a = 8'd76; b = 8'd184;  #10 
a = 8'd76; b = 8'd185;  #10 
a = 8'd76; b = 8'd186;  #10 
a = 8'd76; b = 8'd187;  #10 
a = 8'd76; b = 8'd188;  #10 
a = 8'd76; b = 8'd189;  #10 
a = 8'd76; b = 8'd190;  #10 
a = 8'd76; b = 8'd191;  #10 
a = 8'd76; b = 8'd192;  #10 
a = 8'd76; b = 8'd193;  #10 
a = 8'd76; b = 8'd194;  #10 
a = 8'd76; b = 8'd195;  #10 
a = 8'd76; b = 8'd196;  #10 
a = 8'd76; b = 8'd197;  #10 
a = 8'd76; b = 8'd198;  #10 
a = 8'd76; b = 8'd199;  #10 
a = 8'd76; b = 8'd200;  #10 
a = 8'd76; b = 8'd201;  #10 
a = 8'd76; b = 8'd202;  #10 
a = 8'd76; b = 8'd203;  #10 
a = 8'd76; b = 8'd204;  #10 
a = 8'd76; b = 8'd205;  #10 
a = 8'd76; b = 8'd206;  #10 
a = 8'd76; b = 8'd207;  #10 
a = 8'd76; b = 8'd208;  #10 
a = 8'd76; b = 8'd209;  #10 
a = 8'd76; b = 8'd210;  #10 
a = 8'd76; b = 8'd211;  #10 
a = 8'd76; b = 8'd212;  #10 
a = 8'd76; b = 8'd213;  #10 
a = 8'd76; b = 8'd214;  #10 
a = 8'd76; b = 8'd215;  #10 
a = 8'd76; b = 8'd216;  #10 
a = 8'd76; b = 8'd217;  #10 
a = 8'd76; b = 8'd218;  #10 
a = 8'd76; b = 8'd219;  #10 
a = 8'd76; b = 8'd220;  #10 
a = 8'd76; b = 8'd221;  #10 
a = 8'd76; b = 8'd222;  #10 
a = 8'd76; b = 8'd223;  #10 
a = 8'd76; b = 8'd224;  #10 
a = 8'd76; b = 8'd225;  #10 
a = 8'd76; b = 8'd226;  #10 
a = 8'd76; b = 8'd227;  #10 
a = 8'd76; b = 8'd228;  #10 
a = 8'd76; b = 8'd229;  #10 
a = 8'd76; b = 8'd230;  #10 
a = 8'd76; b = 8'd231;  #10 
a = 8'd76; b = 8'd232;  #10 
a = 8'd76; b = 8'd233;  #10 
a = 8'd76; b = 8'd234;  #10 
a = 8'd76; b = 8'd235;  #10 
a = 8'd76; b = 8'd236;  #10 
a = 8'd76; b = 8'd237;  #10 
a = 8'd76; b = 8'd238;  #10 
a = 8'd76; b = 8'd239;  #10 
a = 8'd76; b = 8'd240;  #10 
a = 8'd76; b = 8'd241;  #10 
a = 8'd76; b = 8'd242;  #10 
a = 8'd76; b = 8'd243;  #10 
a = 8'd76; b = 8'd244;  #10 
a = 8'd76; b = 8'd245;  #10 
a = 8'd76; b = 8'd246;  #10 
a = 8'd76; b = 8'd247;  #10 
a = 8'd76; b = 8'd248;  #10 
a = 8'd76; b = 8'd249;  #10 
a = 8'd76; b = 8'd250;  #10 
a = 8'd76; b = 8'd251;  #10 
a = 8'd76; b = 8'd252;  #10 
a = 8'd76; b = 8'd253;  #10 
a = 8'd76; b = 8'd254;  #10 
a = 8'd76; b = 8'd255;  #10 
a = 8'd77; b = 8'd0;  #10 
a = 8'd77; b = 8'd1;  #10 
a = 8'd77; b = 8'd2;  #10 
a = 8'd77; b = 8'd3;  #10 
a = 8'd77; b = 8'd4;  #10 
a = 8'd77; b = 8'd5;  #10 
a = 8'd77; b = 8'd6;  #10 
a = 8'd77; b = 8'd7;  #10 
a = 8'd77; b = 8'd8;  #10 
a = 8'd77; b = 8'd9;  #10 
a = 8'd77; b = 8'd10;  #10 
a = 8'd77; b = 8'd11;  #10 
a = 8'd77; b = 8'd12;  #10 
a = 8'd77; b = 8'd13;  #10 
a = 8'd77; b = 8'd14;  #10 
a = 8'd77; b = 8'd15;  #10 
a = 8'd77; b = 8'd16;  #10 
a = 8'd77; b = 8'd17;  #10 
a = 8'd77; b = 8'd18;  #10 
a = 8'd77; b = 8'd19;  #10 
a = 8'd77; b = 8'd20;  #10 
a = 8'd77; b = 8'd21;  #10 
a = 8'd77; b = 8'd22;  #10 
a = 8'd77; b = 8'd23;  #10 
a = 8'd77; b = 8'd24;  #10 
a = 8'd77; b = 8'd25;  #10 
a = 8'd77; b = 8'd26;  #10 
a = 8'd77; b = 8'd27;  #10 
a = 8'd77; b = 8'd28;  #10 
a = 8'd77; b = 8'd29;  #10 
a = 8'd77; b = 8'd30;  #10 
a = 8'd77; b = 8'd31;  #10 
a = 8'd77; b = 8'd32;  #10 
a = 8'd77; b = 8'd33;  #10 
a = 8'd77; b = 8'd34;  #10 
a = 8'd77; b = 8'd35;  #10 
a = 8'd77; b = 8'd36;  #10 
a = 8'd77; b = 8'd37;  #10 
a = 8'd77; b = 8'd38;  #10 
a = 8'd77; b = 8'd39;  #10 
a = 8'd77; b = 8'd40;  #10 
a = 8'd77; b = 8'd41;  #10 
a = 8'd77; b = 8'd42;  #10 
a = 8'd77; b = 8'd43;  #10 
a = 8'd77; b = 8'd44;  #10 
a = 8'd77; b = 8'd45;  #10 
a = 8'd77; b = 8'd46;  #10 
a = 8'd77; b = 8'd47;  #10 
a = 8'd77; b = 8'd48;  #10 
a = 8'd77; b = 8'd49;  #10 
a = 8'd77; b = 8'd50;  #10 
a = 8'd77; b = 8'd51;  #10 
a = 8'd77; b = 8'd52;  #10 
a = 8'd77; b = 8'd53;  #10 
a = 8'd77; b = 8'd54;  #10 
a = 8'd77; b = 8'd55;  #10 
a = 8'd77; b = 8'd56;  #10 
a = 8'd77; b = 8'd57;  #10 
a = 8'd77; b = 8'd58;  #10 
a = 8'd77; b = 8'd59;  #10 
a = 8'd77; b = 8'd60;  #10 
a = 8'd77; b = 8'd61;  #10 
a = 8'd77; b = 8'd62;  #10 
a = 8'd77; b = 8'd63;  #10 
a = 8'd77; b = 8'd64;  #10 
a = 8'd77; b = 8'd65;  #10 
a = 8'd77; b = 8'd66;  #10 
a = 8'd77; b = 8'd67;  #10 
a = 8'd77; b = 8'd68;  #10 
a = 8'd77; b = 8'd69;  #10 
a = 8'd77; b = 8'd70;  #10 
a = 8'd77; b = 8'd71;  #10 
a = 8'd77; b = 8'd72;  #10 
a = 8'd77; b = 8'd73;  #10 
a = 8'd77; b = 8'd74;  #10 
a = 8'd77; b = 8'd75;  #10 
a = 8'd77; b = 8'd76;  #10 
a = 8'd77; b = 8'd77;  #10 
a = 8'd77; b = 8'd78;  #10 
a = 8'd77; b = 8'd79;  #10 
a = 8'd77; b = 8'd80;  #10 
a = 8'd77; b = 8'd81;  #10 
a = 8'd77; b = 8'd82;  #10 
a = 8'd77; b = 8'd83;  #10 
a = 8'd77; b = 8'd84;  #10 
a = 8'd77; b = 8'd85;  #10 
a = 8'd77; b = 8'd86;  #10 
a = 8'd77; b = 8'd87;  #10 
a = 8'd77; b = 8'd88;  #10 
a = 8'd77; b = 8'd89;  #10 
a = 8'd77; b = 8'd90;  #10 
a = 8'd77; b = 8'd91;  #10 
a = 8'd77; b = 8'd92;  #10 
a = 8'd77; b = 8'd93;  #10 
a = 8'd77; b = 8'd94;  #10 
a = 8'd77; b = 8'd95;  #10 
a = 8'd77; b = 8'd96;  #10 
a = 8'd77; b = 8'd97;  #10 
a = 8'd77; b = 8'd98;  #10 
a = 8'd77; b = 8'd99;  #10 
a = 8'd77; b = 8'd100;  #10 
a = 8'd77; b = 8'd101;  #10 
a = 8'd77; b = 8'd102;  #10 
a = 8'd77; b = 8'd103;  #10 
a = 8'd77; b = 8'd104;  #10 
a = 8'd77; b = 8'd105;  #10 
a = 8'd77; b = 8'd106;  #10 
a = 8'd77; b = 8'd107;  #10 
a = 8'd77; b = 8'd108;  #10 
a = 8'd77; b = 8'd109;  #10 
a = 8'd77; b = 8'd110;  #10 
a = 8'd77; b = 8'd111;  #10 
a = 8'd77; b = 8'd112;  #10 
a = 8'd77; b = 8'd113;  #10 
a = 8'd77; b = 8'd114;  #10 
a = 8'd77; b = 8'd115;  #10 
a = 8'd77; b = 8'd116;  #10 
a = 8'd77; b = 8'd117;  #10 
a = 8'd77; b = 8'd118;  #10 
a = 8'd77; b = 8'd119;  #10 
a = 8'd77; b = 8'd120;  #10 
a = 8'd77; b = 8'd121;  #10 
a = 8'd77; b = 8'd122;  #10 
a = 8'd77; b = 8'd123;  #10 
a = 8'd77; b = 8'd124;  #10 
a = 8'd77; b = 8'd125;  #10 
a = 8'd77; b = 8'd126;  #10 
a = 8'd77; b = 8'd127;  #10 
a = 8'd77; b = 8'd128;  #10 
a = 8'd77; b = 8'd129;  #10 
a = 8'd77; b = 8'd130;  #10 
a = 8'd77; b = 8'd131;  #10 
a = 8'd77; b = 8'd132;  #10 
a = 8'd77; b = 8'd133;  #10 
a = 8'd77; b = 8'd134;  #10 
a = 8'd77; b = 8'd135;  #10 
a = 8'd77; b = 8'd136;  #10 
a = 8'd77; b = 8'd137;  #10 
a = 8'd77; b = 8'd138;  #10 
a = 8'd77; b = 8'd139;  #10 
a = 8'd77; b = 8'd140;  #10 
a = 8'd77; b = 8'd141;  #10 
a = 8'd77; b = 8'd142;  #10 
a = 8'd77; b = 8'd143;  #10 
a = 8'd77; b = 8'd144;  #10 
a = 8'd77; b = 8'd145;  #10 
a = 8'd77; b = 8'd146;  #10 
a = 8'd77; b = 8'd147;  #10 
a = 8'd77; b = 8'd148;  #10 
a = 8'd77; b = 8'd149;  #10 
a = 8'd77; b = 8'd150;  #10 
a = 8'd77; b = 8'd151;  #10 
a = 8'd77; b = 8'd152;  #10 
a = 8'd77; b = 8'd153;  #10 
a = 8'd77; b = 8'd154;  #10 
a = 8'd77; b = 8'd155;  #10 
a = 8'd77; b = 8'd156;  #10 
a = 8'd77; b = 8'd157;  #10 
a = 8'd77; b = 8'd158;  #10 
a = 8'd77; b = 8'd159;  #10 
a = 8'd77; b = 8'd160;  #10 
a = 8'd77; b = 8'd161;  #10 
a = 8'd77; b = 8'd162;  #10 
a = 8'd77; b = 8'd163;  #10 
a = 8'd77; b = 8'd164;  #10 
a = 8'd77; b = 8'd165;  #10 
a = 8'd77; b = 8'd166;  #10 
a = 8'd77; b = 8'd167;  #10 
a = 8'd77; b = 8'd168;  #10 
a = 8'd77; b = 8'd169;  #10 
a = 8'd77; b = 8'd170;  #10 
a = 8'd77; b = 8'd171;  #10 
a = 8'd77; b = 8'd172;  #10 
a = 8'd77; b = 8'd173;  #10 
a = 8'd77; b = 8'd174;  #10 
a = 8'd77; b = 8'd175;  #10 
a = 8'd77; b = 8'd176;  #10 
a = 8'd77; b = 8'd177;  #10 
a = 8'd77; b = 8'd178;  #10 
a = 8'd77; b = 8'd179;  #10 
a = 8'd77; b = 8'd180;  #10 
a = 8'd77; b = 8'd181;  #10 
a = 8'd77; b = 8'd182;  #10 
a = 8'd77; b = 8'd183;  #10 
a = 8'd77; b = 8'd184;  #10 
a = 8'd77; b = 8'd185;  #10 
a = 8'd77; b = 8'd186;  #10 
a = 8'd77; b = 8'd187;  #10 
a = 8'd77; b = 8'd188;  #10 
a = 8'd77; b = 8'd189;  #10 
a = 8'd77; b = 8'd190;  #10 
a = 8'd77; b = 8'd191;  #10 
a = 8'd77; b = 8'd192;  #10 
a = 8'd77; b = 8'd193;  #10 
a = 8'd77; b = 8'd194;  #10 
a = 8'd77; b = 8'd195;  #10 
a = 8'd77; b = 8'd196;  #10 
a = 8'd77; b = 8'd197;  #10 
a = 8'd77; b = 8'd198;  #10 
a = 8'd77; b = 8'd199;  #10 
a = 8'd77; b = 8'd200;  #10 
a = 8'd77; b = 8'd201;  #10 
a = 8'd77; b = 8'd202;  #10 
a = 8'd77; b = 8'd203;  #10 
a = 8'd77; b = 8'd204;  #10 
a = 8'd77; b = 8'd205;  #10 
a = 8'd77; b = 8'd206;  #10 
a = 8'd77; b = 8'd207;  #10 
a = 8'd77; b = 8'd208;  #10 
a = 8'd77; b = 8'd209;  #10 
a = 8'd77; b = 8'd210;  #10 
a = 8'd77; b = 8'd211;  #10 
a = 8'd77; b = 8'd212;  #10 
a = 8'd77; b = 8'd213;  #10 
a = 8'd77; b = 8'd214;  #10 
a = 8'd77; b = 8'd215;  #10 
a = 8'd77; b = 8'd216;  #10 
a = 8'd77; b = 8'd217;  #10 
a = 8'd77; b = 8'd218;  #10 
a = 8'd77; b = 8'd219;  #10 
a = 8'd77; b = 8'd220;  #10 
a = 8'd77; b = 8'd221;  #10 
a = 8'd77; b = 8'd222;  #10 
a = 8'd77; b = 8'd223;  #10 
a = 8'd77; b = 8'd224;  #10 
a = 8'd77; b = 8'd225;  #10 
a = 8'd77; b = 8'd226;  #10 
a = 8'd77; b = 8'd227;  #10 
a = 8'd77; b = 8'd228;  #10 
a = 8'd77; b = 8'd229;  #10 
a = 8'd77; b = 8'd230;  #10 
a = 8'd77; b = 8'd231;  #10 
a = 8'd77; b = 8'd232;  #10 
a = 8'd77; b = 8'd233;  #10 
a = 8'd77; b = 8'd234;  #10 
a = 8'd77; b = 8'd235;  #10 
a = 8'd77; b = 8'd236;  #10 
a = 8'd77; b = 8'd237;  #10 
a = 8'd77; b = 8'd238;  #10 
a = 8'd77; b = 8'd239;  #10 
a = 8'd77; b = 8'd240;  #10 
a = 8'd77; b = 8'd241;  #10 
a = 8'd77; b = 8'd242;  #10 
a = 8'd77; b = 8'd243;  #10 
a = 8'd77; b = 8'd244;  #10 
a = 8'd77; b = 8'd245;  #10 
a = 8'd77; b = 8'd246;  #10 
a = 8'd77; b = 8'd247;  #10 
a = 8'd77; b = 8'd248;  #10 
a = 8'd77; b = 8'd249;  #10 
a = 8'd77; b = 8'd250;  #10 
a = 8'd77; b = 8'd251;  #10 
a = 8'd77; b = 8'd252;  #10 
a = 8'd77; b = 8'd253;  #10 
a = 8'd77; b = 8'd254;  #10 
a = 8'd77; b = 8'd255;  #10 
a = 8'd78; b = 8'd0;  #10 
a = 8'd78; b = 8'd1;  #10 
a = 8'd78; b = 8'd2;  #10 
a = 8'd78; b = 8'd3;  #10 
a = 8'd78; b = 8'd4;  #10 
a = 8'd78; b = 8'd5;  #10 
a = 8'd78; b = 8'd6;  #10 
a = 8'd78; b = 8'd7;  #10 
a = 8'd78; b = 8'd8;  #10 
a = 8'd78; b = 8'd9;  #10 
a = 8'd78; b = 8'd10;  #10 
a = 8'd78; b = 8'd11;  #10 
a = 8'd78; b = 8'd12;  #10 
a = 8'd78; b = 8'd13;  #10 
a = 8'd78; b = 8'd14;  #10 
a = 8'd78; b = 8'd15;  #10 
a = 8'd78; b = 8'd16;  #10 
a = 8'd78; b = 8'd17;  #10 
a = 8'd78; b = 8'd18;  #10 
a = 8'd78; b = 8'd19;  #10 
a = 8'd78; b = 8'd20;  #10 
a = 8'd78; b = 8'd21;  #10 
a = 8'd78; b = 8'd22;  #10 
a = 8'd78; b = 8'd23;  #10 
a = 8'd78; b = 8'd24;  #10 
a = 8'd78; b = 8'd25;  #10 
a = 8'd78; b = 8'd26;  #10 
a = 8'd78; b = 8'd27;  #10 
a = 8'd78; b = 8'd28;  #10 
a = 8'd78; b = 8'd29;  #10 
a = 8'd78; b = 8'd30;  #10 
a = 8'd78; b = 8'd31;  #10 
a = 8'd78; b = 8'd32;  #10 
a = 8'd78; b = 8'd33;  #10 
a = 8'd78; b = 8'd34;  #10 
a = 8'd78; b = 8'd35;  #10 
a = 8'd78; b = 8'd36;  #10 
a = 8'd78; b = 8'd37;  #10 
a = 8'd78; b = 8'd38;  #10 
a = 8'd78; b = 8'd39;  #10 
a = 8'd78; b = 8'd40;  #10 
a = 8'd78; b = 8'd41;  #10 
a = 8'd78; b = 8'd42;  #10 
a = 8'd78; b = 8'd43;  #10 
a = 8'd78; b = 8'd44;  #10 
a = 8'd78; b = 8'd45;  #10 
a = 8'd78; b = 8'd46;  #10 
a = 8'd78; b = 8'd47;  #10 
a = 8'd78; b = 8'd48;  #10 
a = 8'd78; b = 8'd49;  #10 
a = 8'd78; b = 8'd50;  #10 
a = 8'd78; b = 8'd51;  #10 
a = 8'd78; b = 8'd52;  #10 
a = 8'd78; b = 8'd53;  #10 
a = 8'd78; b = 8'd54;  #10 
a = 8'd78; b = 8'd55;  #10 
a = 8'd78; b = 8'd56;  #10 
a = 8'd78; b = 8'd57;  #10 
a = 8'd78; b = 8'd58;  #10 
a = 8'd78; b = 8'd59;  #10 
a = 8'd78; b = 8'd60;  #10 
a = 8'd78; b = 8'd61;  #10 
a = 8'd78; b = 8'd62;  #10 
a = 8'd78; b = 8'd63;  #10 
a = 8'd78; b = 8'd64;  #10 
a = 8'd78; b = 8'd65;  #10 
a = 8'd78; b = 8'd66;  #10 
a = 8'd78; b = 8'd67;  #10 
a = 8'd78; b = 8'd68;  #10 
a = 8'd78; b = 8'd69;  #10 
a = 8'd78; b = 8'd70;  #10 
a = 8'd78; b = 8'd71;  #10 
a = 8'd78; b = 8'd72;  #10 
a = 8'd78; b = 8'd73;  #10 
a = 8'd78; b = 8'd74;  #10 
a = 8'd78; b = 8'd75;  #10 
a = 8'd78; b = 8'd76;  #10 
a = 8'd78; b = 8'd77;  #10 
a = 8'd78; b = 8'd78;  #10 
a = 8'd78; b = 8'd79;  #10 
a = 8'd78; b = 8'd80;  #10 
a = 8'd78; b = 8'd81;  #10 
a = 8'd78; b = 8'd82;  #10 
a = 8'd78; b = 8'd83;  #10 
a = 8'd78; b = 8'd84;  #10 
a = 8'd78; b = 8'd85;  #10 
a = 8'd78; b = 8'd86;  #10 
a = 8'd78; b = 8'd87;  #10 
a = 8'd78; b = 8'd88;  #10 
a = 8'd78; b = 8'd89;  #10 
a = 8'd78; b = 8'd90;  #10 
a = 8'd78; b = 8'd91;  #10 
a = 8'd78; b = 8'd92;  #10 
a = 8'd78; b = 8'd93;  #10 
a = 8'd78; b = 8'd94;  #10 
a = 8'd78; b = 8'd95;  #10 
a = 8'd78; b = 8'd96;  #10 
a = 8'd78; b = 8'd97;  #10 
a = 8'd78; b = 8'd98;  #10 
a = 8'd78; b = 8'd99;  #10 
a = 8'd78; b = 8'd100;  #10 
a = 8'd78; b = 8'd101;  #10 
a = 8'd78; b = 8'd102;  #10 
a = 8'd78; b = 8'd103;  #10 
a = 8'd78; b = 8'd104;  #10 
a = 8'd78; b = 8'd105;  #10 
a = 8'd78; b = 8'd106;  #10 
a = 8'd78; b = 8'd107;  #10 
a = 8'd78; b = 8'd108;  #10 
a = 8'd78; b = 8'd109;  #10 
a = 8'd78; b = 8'd110;  #10 
a = 8'd78; b = 8'd111;  #10 
a = 8'd78; b = 8'd112;  #10 
a = 8'd78; b = 8'd113;  #10 
a = 8'd78; b = 8'd114;  #10 
a = 8'd78; b = 8'd115;  #10 
a = 8'd78; b = 8'd116;  #10 
a = 8'd78; b = 8'd117;  #10 
a = 8'd78; b = 8'd118;  #10 
a = 8'd78; b = 8'd119;  #10 
a = 8'd78; b = 8'd120;  #10 
a = 8'd78; b = 8'd121;  #10 
a = 8'd78; b = 8'd122;  #10 
a = 8'd78; b = 8'd123;  #10 
a = 8'd78; b = 8'd124;  #10 
a = 8'd78; b = 8'd125;  #10 
a = 8'd78; b = 8'd126;  #10 
a = 8'd78; b = 8'd127;  #10 
a = 8'd78; b = 8'd128;  #10 
a = 8'd78; b = 8'd129;  #10 
a = 8'd78; b = 8'd130;  #10 
a = 8'd78; b = 8'd131;  #10 
a = 8'd78; b = 8'd132;  #10 
a = 8'd78; b = 8'd133;  #10 
a = 8'd78; b = 8'd134;  #10 
a = 8'd78; b = 8'd135;  #10 
a = 8'd78; b = 8'd136;  #10 
a = 8'd78; b = 8'd137;  #10 
a = 8'd78; b = 8'd138;  #10 
a = 8'd78; b = 8'd139;  #10 
a = 8'd78; b = 8'd140;  #10 
a = 8'd78; b = 8'd141;  #10 
a = 8'd78; b = 8'd142;  #10 
a = 8'd78; b = 8'd143;  #10 
a = 8'd78; b = 8'd144;  #10 
a = 8'd78; b = 8'd145;  #10 
a = 8'd78; b = 8'd146;  #10 
a = 8'd78; b = 8'd147;  #10 
a = 8'd78; b = 8'd148;  #10 
a = 8'd78; b = 8'd149;  #10 
a = 8'd78; b = 8'd150;  #10 
a = 8'd78; b = 8'd151;  #10 
a = 8'd78; b = 8'd152;  #10 
a = 8'd78; b = 8'd153;  #10 
a = 8'd78; b = 8'd154;  #10 
a = 8'd78; b = 8'd155;  #10 
a = 8'd78; b = 8'd156;  #10 
a = 8'd78; b = 8'd157;  #10 
a = 8'd78; b = 8'd158;  #10 
a = 8'd78; b = 8'd159;  #10 
a = 8'd78; b = 8'd160;  #10 
a = 8'd78; b = 8'd161;  #10 
a = 8'd78; b = 8'd162;  #10 
a = 8'd78; b = 8'd163;  #10 
a = 8'd78; b = 8'd164;  #10 
a = 8'd78; b = 8'd165;  #10 
a = 8'd78; b = 8'd166;  #10 
a = 8'd78; b = 8'd167;  #10 
a = 8'd78; b = 8'd168;  #10 
a = 8'd78; b = 8'd169;  #10 
a = 8'd78; b = 8'd170;  #10 
a = 8'd78; b = 8'd171;  #10 
a = 8'd78; b = 8'd172;  #10 
a = 8'd78; b = 8'd173;  #10 
a = 8'd78; b = 8'd174;  #10 
a = 8'd78; b = 8'd175;  #10 
a = 8'd78; b = 8'd176;  #10 
a = 8'd78; b = 8'd177;  #10 
a = 8'd78; b = 8'd178;  #10 
a = 8'd78; b = 8'd179;  #10 
a = 8'd78; b = 8'd180;  #10 
a = 8'd78; b = 8'd181;  #10 
a = 8'd78; b = 8'd182;  #10 
a = 8'd78; b = 8'd183;  #10 
a = 8'd78; b = 8'd184;  #10 
a = 8'd78; b = 8'd185;  #10 
a = 8'd78; b = 8'd186;  #10 
a = 8'd78; b = 8'd187;  #10 
a = 8'd78; b = 8'd188;  #10 
a = 8'd78; b = 8'd189;  #10 
a = 8'd78; b = 8'd190;  #10 
a = 8'd78; b = 8'd191;  #10 
a = 8'd78; b = 8'd192;  #10 
a = 8'd78; b = 8'd193;  #10 
a = 8'd78; b = 8'd194;  #10 
a = 8'd78; b = 8'd195;  #10 
a = 8'd78; b = 8'd196;  #10 
a = 8'd78; b = 8'd197;  #10 
a = 8'd78; b = 8'd198;  #10 
a = 8'd78; b = 8'd199;  #10 
a = 8'd78; b = 8'd200;  #10 
a = 8'd78; b = 8'd201;  #10 
a = 8'd78; b = 8'd202;  #10 
a = 8'd78; b = 8'd203;  #10 
a = 8'd78; b = 8'd204;  #10 
a = 8'd78; b = 8'd205;  #10 
a = 8'd78; b = 8'd206;  #10 
a = 8'd78; b = 8'd207;  #10 
a = 8'd78; b = 8'd208;  #10 
a = 8'd78; b = 8'd209;  #10 
a = 8'd78; b = 8'd210;  #10 
a = 8'd78; b = 8'd211;  #10 
a = 8'd78; b = 8'd212;  #10 
a = 8'd78; b = 8'd213;  #10 
a = 8'd78; b = 8'd214;  #10 
a = 8'd78; b = 8'd215;  #10 
a = 8'd78; b = 8'd216;  #10 
a = 8'd78; b = 8'd217;  #10 
a = 8'd78; b = 8'd218;  #10 
a = 8'd78; b = 8'd219;  #10 
a = 8'd78; b = 8'd220;  #10 
a = 8'd78; b = 8'd221;  #10 
a = 8'd78; b = 8'd222;  #10 
a = 8'd78; b = 8'd223;  #10 
a = 8'd78; b = 8'd224;  #10 
a = 8'd78; b = 8'd225;  #10 
a = 8'd78; b = 8'd226;  #10 
a = 8'd78; b = 8'd227;  #10 
a = 8'd78; b = 8'd228;  #10 
a = 8'd78; b = 8'd229;  #10 
a = 8'd78; b = 8'd230;  #10 
a = 8'd78; b = 8'd231;  #10 
a = 8'd78; b = 8'd232;  #10 
a = 8'd78; b = 8'd233;  #10 
a = 8'd78; b = 8'd234;  #10 
a = 8'd78; b = 8'd235;  #10 
a = 8'd78; b = 8'd236;  #10 
a = 8'd78; b = 8'd237;  #10 
a = 8'd78; b = 8'd238;  #10 
a = 8'd78; b = 8'd239;  #10 
a = 8'd78; b = 8'd240;  #10 
a = 8'd78; b = 8'd241;  #10 
a = 8'd78; b = 8'd242;  #10 
a = 8'd78; b = 8'd243;  #10 
a = 8'd78; b = 8'd244;  #10 
a = 8'd78; b = 8'd245;  #10 
a = 8'd78; b = 8'd246;  #10 
a = 8'd78; b = 8'd247;  #10 
a = 8'd78; b = 8'd248;  #10 
a = 8'd78; b = 8'd249;  #10 
a = 8'd78; b = 8'd250;  #10 
a = 8'd78; b = 8'd251;  #10 
a = 8'd78; b = 8'd252;  #10 
a = 8'd78; b = 8'd253;  #10 
a = 8'd78; b = 8'd254;  #10 
a = 8'd78; b = 8'd255;  #10 
a = 8'd79; b = 8'd0;  #10 
a = 8'd79; b = 8'd1;  #10 
a = 8'd79; b = 8'd2;  #10 
a = 8'd79; b = 8'd3;  #10 
a = 8'd79; b = 8'd4;  #10 
a = 8'd79; b = 8'd5;  #10 
a = 8'd79; b = 8'd6;  #10 
a = 8'd79; b = 8'd7;  #10 
a = 8'd79; b = 8'd8;  #10 
a = 8'd79; b = 8'd9;  #10 
a = 8'd79; b = 8'd10;  #10 
a = 8'd79; b = 8'd11;  #10 
a = 8'd79; b = 8'd12;  #10 
a = 8'd79; b = 8'd13;  #10 
a = 8'd79; b = 8'd14;  #10 
a = 8'd79; b = 8'd15;  #10 
a = 8'd79; b = 8'd16;  #10 
a = 8'd79; b = 8'd17;  #10 
a = 8'd79; b = 8'd18;  #10 
a = 8'd79; b = 8'd19;  #10 
a = 8'd79; b = 8'd20;  #10 
a = 8'd79; b = 8'd21;  #10 
a = 8'd79; b = 8'd22;  #10 
a = 8'd79; b = 8'd23;  #10 
a = 8'd79; b = 8'd24;  #10 
a = 8'd79; b = 8'd25;  #10 
a = 8'd79; b = 8'd26;  #10 
a = 8'd79; b = 8'd27;  #10 
a = 8'd79; b = 8'd28;  #10 
a = 8'd79; b = 8'd29;  #10 
a = 8'd79; b = 8'd30;  #10 
a = 8'd79; b = 8'd31;  #10 
a = 8'd79; b = 8'd32;  #10 
a = 8'd79; b = 8'd33;  #10 
a = 8'd79; b = 8'd34;  #10 
a = 8'd79; b = 8'd35;  #10 
a = 8'd79; b = 8'd36;  #10 
a = 8'd79; b = 8'd37;  #10 
a = 8'd79; b = 8'd38;  #10 
a = 8'd79; b = 8'd39;  #10 
a = 8'd79; b = 8'd40;  #10 
a = 8'd79; b = 8'd41;  #10 
a = 8'd79; b = 8'd42;  #10 
a = 8'd79; b = 8'd43;  #10 
a = 8'd79; b = 8'd44;  #10 
a = 8'd79; b = 8'd45;  #10 
a = 8'd79; b = 8'd46;  #10 
a = 8'd79; b = 8'd47;  #10 
a = 8'd79; b = 8'd48;  #10 
a = 8'd79; b = 8'd49;  #10 
a = 8'd79; b = 8'd50;  #10 
a = 8'd79; b = 8'd51;  #10 
a = 8'd79; b = 8'd52;  #10 
a = 8'd79; b = 8'd53;  #10 
a = 8'd79; b = 8'd54;  #10 
a = 8'd79; b = 8'd55;  #10 
a = 8'd79; b = 8'd56;  #10 
a = 8'd79; b = 8'd57;  #10 
a = 8'd79; b = 8'd58;  #10 
a = 8'd79; b = 8'd59;  #10 
a = 8'd79; b = 8'd60;  #10 
a = 8'd79; b = 8'd61;  #10 
a = 8'd79; b = 8'd62;  #10 
a = 8'd79; b = 8'd63;  #10 
a = 8'd79; b = 8'd64;  #10 
a = 8'd79; b = 8'd65;  #10 
a = 8'd79; b = 8'd66;  #10 
a = 8'd79; b = 8'd67;  #10 
a = 8'd79; b = 8'd68;  #10 
a = 8'd79; b = 8'd69;  #10 
a = 8'd79; b = 8'd70;  #10 
a = 8'd79; b = 8'd71;  #10 
a = 8'd79; b = 8'd72;  #10 
a = 8'd79; b = 8'd73;  #10 
a = 8'd79; b = 8'd74;  #10 
a = 8'd79; b = 8'd75;  #10 
a = 8'd79; b = 8'd76;  #10 
a = 8'd79; b = 8'd77;  #10 
a = 8'd79; b = 8'd78;  #10 
a = 8'd79; b = 8'd79;  #10 
a = 8'd79; b = 8'd80;  #10 
a = 8'd79; b = 8'd81;  #10 
a = 8'd79; b = 8'd82;  #10 
a = 8'd79; b = 8'd83;  #10 
a = 8'd79; b = 8'd84;  #10 
a = 8'd79; b = 8'd85;  #10 
a = 8'd79; b = 8'd86;  #10 
a = 8'd79; b = 8'd87;  #10 
a = 8'd79; b = 8'd88;  #10 
a = 8'd79; b = 8'd89;  #10 
a = 8'd79; b = 8'd90;  #10 
a = 8'd79; b = 8'd91;  #10 
a = 8'd79; b = 8'd92;  #10 
a = 8'd79; b = 8'd93;  #10 
a = 8'd79; b = 8'd94;  #10 
a = 8'd79; b = 8'd95;  #10 
a = 8'd79; b = 8'd96;  #10 
a = 8'd79; b = 8'd97;  #10 
a = 8'd79; b = 8'd98;  #10 
a = 8'd79; b = 8'd99;  #10 
a = 8'd79; b = 8'd100;  #10 
a = 8'd79; b = 8'd101;  #10 
a = 8'd79; b = 8'd102;  #10 
a = 8'd79; b = 8'd103;  #10 
a = 8'd79; b = 8'd104;  #10 
a = 8'd79; b = 8'd105;  #10 
a = 8'd79; b = 8'd106;  #10 
a = 8'd79; b = 8'd107;  #10 
a = 8'd79; b = 8'd108;  #10 
a = 8'd79; b = 8'd109;  #10 
a = 8'd79; b = 8'd110;  #10 
a = 8'd79; b = 8'd111;  #10 
a = 8'd79; b = 8'd112;  #10 
a = 8'd79; b = 8'd113;  #10 
a = 8'd79; b = 8'd114;  #10 
a = 8'd79; b = 8'd115;  #10 
a = 8'd79; b = 8'd116;  #10 
a = 8'd79; b = 8'd117;  #10 
a = 8'd79; b = 8'd118;  #10 
a = 8'd79; b = 8'd119;  #10 
a = 8'd79; b = 8'd120;  #10 
a = 8'd79; b = 8'd121;  #10 
a = 8'd79; b = 8'd122;  #10 
a = 8'd79; b = 8'd123;  #10 
a = 8'd79; b = 8'd124;  #10 
a = 8'd79; b = 8'd125;  #10 
a = 8'd79; b = 8'd126;  #10 
a = 8'd79; b = 8'd127;  #10 
a = 8'd79; b = 8'd128;  #10 
a = 8'd79; b = 8'd129;  #10 
a = 8'd79; b = 8'd130;  #10 
a = 8'd79; b = 8'd131;  #10 
a = 8'd79; b = 8'd132;  #10 
a = 8'd79; b = 8'd133;  #10 
a = 8'd79; b = 8'd134;  #10 
a = 8'd79; b = 8'd135;  #10 
a = 8'd79; b = 8'd136;  #10 
a = 8'd79; b = 8'd137;  #10 
a = 8'd79; b = 8'd138;  #10 
a = 8'd79; b = 8'd139;  #10 
a = 8'd79; b = 8'd140;  #10 
a = 8'd79; b = 8'd141;  #10 
a = 8'd79; b = 8'd142;  #10 
a = 8'd79; b = 8'd143;  #10 
a = 8'd79; b = 8'd144;  #10 
a = 8'd79; b = 8'd145;  #10 
a = 8'd79; b = 8'd146;  #10 
a = 8'd79; b = 8'd147;  #10 
a = 8'd79; b = 8'd148;  #10 
a = 8'd79; b = 8'd149;  #10 
a = 8'd79; b = 8'd150;  #10 
a = 8'd79; b = 8'd151;  #10 
a = 8'd79; b = 8'd152;  #10 
a = 8'd79; b = 8'd153;  #10 
a = 8'd79; b = 8'd154;  #10 
a = 8'd79; b = 8'd155;  #10 
a = 8'd79; b = 8'd156;  #10 
a = 8'd79; b = 8'd157;  #10 
a = 8'd79; b = 8'd158;  #10 
a = 8'd79; b = 8'd159;  #10 
a = 8'd79; b = 8'd160;  #10 
a = 8'd79; b = 8'd161;  #10 
a = 8'd79; b = 8'd162;  #10 
a = 8'd79; b = 8'd163;  #10 
a = 8'd79; b = 8'd164;  #10 
a = 8'd79; b = 8'd165;  #10 
a = 8'd79; b = 8'd166;  #10 
a = 8'd79; b = 8'd167;  #10 
a = 8'd79; b = 8'd168;  #10 
a = 8'd79; b = 8'd169;  #10 
a = 8'd79; b = 8'd170;  #10 
a = 8'd79; b = 8'd171;  #10 
a = 8'd79; b = 8'd172;  #10 
a = 8'd79; b = 8'd173;  #10 
a = 8'd79; b = 8'd174;  #10 
a = 8'd79; b = 8'd175;  #10 
a = 8'd79; b = 8'd176;  #10 
a = 8'd79; b = 8'd177;  #10 
a = 8'd79; b = 8'd178;  #10 
a = 8'd79; b = 8'd179;  #10 
a = 8'd79; b = 8'd180;  #10 
a = 8'd79; b = 8'd181;  #10 
a = 8'd79; b = 8'd182;  #10 
a = 8'd79; b = 8'd183;  #10 
a = 8'd79; b = 8'd184;  #10 
a = 8'd79; b = 8'd185;  #10 
a = 8'd79; b = 8'd186;  #10 
a = 8'd79; b = 8'd187;  #10 
a = 8'd79; b = 8'd188;  #10 
a = 8'd79; b = 8'd189;  #10 
a = 8'd79; b = 8'd190;  #10 
a = 8'd79; b = 8'd191;  #10 
a = 8'd79; b = 8'd192;  #10 
a = 8'd79; b = 8'd193;  #10 
a = 8'd79; b = 8'd194;  #10 
a = 8'd79; b = 8'd195;  #10 
a = 8'd79; b = 8'd196;  #10 
a = 8'd79; b = 8'd197;  #10 
a = 8'd79; b = 8'd198;  #10 
a = 8'd79; b = 8'd199;  #10 
a = 8'd79; b = 8'd200;  #10 
a = 8'd79; b = 8'd201;  #10 
a = 8'd79; b = 8'd202;  #10 
a = 8'd79; b = 8'd203;  #10 
a = 8'd79; b = 8'd204;  #10 
a = 8'd79; b = 8'd205;  #10 
a = 8'd79; b = 8'd206;  #10 
a = 8'd79; b = 8'd207;  #10 
a = 8'd79; b = 8'd208;  #10 
a = 8'd79; b = 8'd209;  #10 
a = 8'd79; b = 8'd210;  #10 
a = 8'd79; b = 8'd211;  #10 
a = 8'd79; b = 8'd212;  #10 
a = 8'd79; b = 8'd213;  #10 
a = 8'd79; b = 8'd214;  #10 
a = 8'd79; b = 8'd215;  #10 
a = 8'd79; b = 8'd216;  #10 
a = 8'd79; b = 8'd217;  #10 
a = 8'd79; b = 8'd218;  #10 
a = 8'd79; b = 8'd219;  #10 
a = 8'd79; b = 8'd220;  #10 
a = 8'd79; b = 8'd221;  #10 
a = 8'd79; b = 8'd222;  #10 
a = 8'd79; b = 8'd223;  #10 
a = 8'd79; b = 8'd224;  #10 
a = 8'd79; b = 8'd225;  #10 
a = 8'd79; b = 8'd226;  #10 
a = 8'd79; b = 8'd227;  #10 
a = 8'd79; b = 8'd228;  #10 
a = 8'd79; b = 8'd229;  #10 
a = 8'd79; b = 8'd230;  #10 
a = 8'd79; b = 8'd231;  #10 
a = 8'd79; b = 8'd232;  #10 
a = 8'd79; b = 8'd233;  #10 
a = 8'd79; b = 8'd234;  #10 
a = 8'd79; b = 8'd235;  #10 
a = 8'd79; b = 8'd236;  #10 
a = 8'd79; b = 8'd237;  #10 
a = 8'd79; b = 8'd238;  #10 
a = 8'd79; b = 8'd239;  #10 
a = 8'd79; b = 8'd240;  #10 
a = 8'd79; b = 8'd241;  #10 
a = 8'd79; b = 8'd242;  #10 
a = 8'd79; b = 8'd243;  #10 
a = 8'd79; b = 8'd244;  #10 
a = 8'd79; b = 8'd245;  #10 
a = 8'd79; b = 8'd246;  #10 
a = 8'd79; b = 8'd247;  #10 
a = 8'd79; b = 8'd248;  #10 
a = 8'd79; b = 8'd249;  #10 
a = 8'd79; b = 8'd250;  #10 
a = 8'd79; b = 8'd251;  #10 
a = 8'd79; b = 8'd252;  #10 
a = 8'd79; b = 8'd253;  #10 
a = 8'd79; b = 8'd254;  #10 
a = 8'd79; b = 8'd255;  #10 
a = 8'd80; b = 8'd0;  #10 
a = 8'd80; b = 8'd1;  #10 
a = 8'd80; b = 8'd2;  #10 
a = 8'd80; b = 8'd3;  #10 
a = 8'd80; b = 8'd4;  #10 
a = 8'd80; b = 8'd5;  #10 
a = 8'd80; b = 8'd6;  #10 
a = 8'd80; b = 8'd7;  #10 
a = 8'd80; b = 8'd8;  #10 
a = 8'd80; b = 8'd9;  #10 
a = 8'd80; b = 8'd10;  #10 
a = 8'd80; b = 8'd11;  #10 
a = 8'd80; b = 8'd12;  #10 
a = 8'd80; b = 8'd13;  #10 
a = 8'd80; b = 8'd14;  #10 
a = 8'd80; b = 8'd15;  #10 
a = 8'd80; b = 8'd16;  #10 
a = 8'd80; b = 8'd17;  #10 
a = 8'd80; b = 8'd18;  #10 
a = 8'd80; b = 8'd19;  #10 
a = 8'd80; b = 8'd20;  #10 
a = 8'd80; b = 8'd21;  #10 
a = 8'd80; b = 8'd22;  #10 
a = 8'd80; b = 8'd23;  #10 
a = 8'd80; b = 8'd24;  #10 
a = 8'd80; b = 8'd25;  #10 
a = 8'd80; b = 8'd26;  #10 
a = 8'd80; b = 8'd27;  #10 
a = 8'd80; b = 8'd28;  #10 
a = 8'd80; b = 8'd29;  #10 
a = 8'd80; b = 8'd30;  #10 
a = 8'd80; b = 8'd31;  #10 
a = 8'd80; b = 8'd32;  #10 
a = 8'd80; b = 8'd33;  #10 
a = 8'd80; b = 8'd34;  #10 
a = 8'd80; b = 8'd35;  #10 
a = 8'd80; b = 8'd36;  #10 
a = 8'd80; b = 8'd37;  #10 
a = 8'd80; b = 8'd38;  #10 
a = 8'd80; b = 8'd39;  #10 
a = 8'd80; b = 8'd40;  #10 
a = 8'd80; b = 8'd41;  #10 
a = 8'd80; b = 8'd42;  #10 
a = 8'd80; b = 8'd43;  #10 
a = 8'd80; b = 8'd44;  #10 
a = 8'd80; b = 8'd45;  #10 
a = 8'd80; b = 8'd46;  #10 
a = 8'd80; b = 8'd47;  #10 
a = 8'd80; b = 8'd48;  #10 
a = 8'd80; b = 8'd49;  #10 
a = 8'd80; b = 8'd50;  #10 
a = 8'd80; b = 8'd51;  #10 
a = 8'd80; b = 8'd52;  #10 
a = 8'd80; b = 8'd53;  #10 
a = 8'd80; b = 8'd54;  #10 
a = 8'd80; b = 8'd55;  #10 
a = 8'd80; b = 8'd56;  #10 
a = 8'd80; b = 8'd57;  #10 
a = 8'd80; b = 8'd58;  #10 
a = 8'd80; b = 8'd59;  #10 
a = 8'd80; b = 8'd60;  #10 
a = 8'd80; b = 8'd61;  #10 
a = 8'd80; b = 8'd62;  #10 
a = 8'd80; b = 8'd63;  #10 
a = 8'd80; b = 8'd64;  #10 
a = 8'd80; b = 8'd65;  #10 
a = 8'd80; b = 8'd66;  #10 
a = 8'd80; b = 8'd67;  #10 
a = 8'd80; b = 8'd68;  #10 
a = 8'd80; b = 8'd69;  #10 
a = 8'd80; b = 8'd70;  #10 
a = 8'd80; b = 8'd71;  #10 
a = 8'd80; b = 8'd72;  #10 
a = 8'd80; b = 8'd73;  #10 
a = 8'd80; b = 8'd74;  #10 
a = 8'd80; b = 8'd75;  #10 
a = 8'd80; b = 8'd76;  #10 
a = 8'd80; b = 8'd77;  #10 
a = 8'd80; b = 8'd78;  #10 
a = 8'd80; b = 8'd79;  #10 
a = 8'd80; b = 8'd80;  #10 
a = 8'd80; b = 8'd81;  #10 
a = 8'd80; b = 8'd82;  #10 
a = 8'd80; b = 8'd83;  #10 
a = 8'd80; b = 8'd84;  #10 
a = 8'd80; b = 8'd85;  #10 
a = 8'd80; b = 8'd86;  #10 
a = 8'd80; b = 8'd87;  #10 
a = 8'd80; b = 8'd88;  #10 
a = 8'd80; b = 8'd89;  #10 
a = 8'd80; b = 8'd90;  #10 
a = 8'd80; b = 8'd91;  #10 
a = 8'd80; b = 8'd92;  #10 
a = 8'd80; b = 8'd93;  #10 
a = 8'd80; b = 8'd94;  #10 
a = 8'd80; b = 8'd95;  #10 
a = 8'd80; b = 8'd96;  #10 
a = 8'd80; b = 8'd97;  #10 
a = 8'd80; b = 8'd98;  #10 
a = 8'd80; b = 8'd99;  #10 
a = 8'd80; b = 8'd100;  #10 
a = 8'd80; b = 8'd101;  #10 
a = 8'd80; b = 8'd102;  #10 
a = 8'd80; b = 8'd103;  #10 
a = 8'd80; b = 8'd104;  #10 
a = 8'd80; b = 8'd105;  #10 
a = 8'd80; b = 8'd106;  #10 
a = 8'd80; b = 8'd107;  #10 
a = 8'd80; b = 8'd108;  #10 
a = 8'd80; b = 8'd109;  #10 
a = 8'd80; b = 8'd110;  #10 
a = 8'd80; b = 8'd111;  #10 
a = 8'd80; b = 8'd112;  #10 
a = 8'd80; b = 8'd113;  #10 
a = 8'd80; b = 8'd114;  #10 
a = 8'd80; b = 8'd115;  #10 
a = 8'd80; b = 8'd116;  #10 
a = 8'd80; b = 8'd117;  #10 
a = 8'd80; b = 8'd118;  #10 
a = 8'd80; b = 8'd119;  #10 
a = 8'd80; b = 8'd120;  #10 
a = 8'd80; b = 8'd121;  #10 
a = 8'd80; b = 8'd122;  #10 
a = 8'd80; b = 8'd123;  #10 
a = 8'd80; b = 8'd124;  #10 
a = 8'd80; b = 8'd125;  #10 
a = 8'd80; b = 8'd126;  #10 
a = 8'd80; b = 8'd127;  #10 
a = 8'd80; b = 8'd128;  #10 
a = 8'd80; b = 8'd129;  #10 
a = 8'd80; b = 8'd130;  #10 
a = 8'd80; b = 8'd131;  #10 
a = 8'd80; b = 8'd132;  #10 
a = 8'd80; b = 8'd133;  #10 
a = 8'd80; b = 8'd134;  #10 
a = 8'd80; b = 8'd135;  #10 
a = 8'd80; b = 8'd136;  #10 
a = 8'd80; b = 8'd137;  #10 
a = 8'd80; b = 8'd138;  #10 
a = 8'd80; b = 8'd139;  #10 
a = 8'd80; b = 8'd140;  #10 
a = 8'd80; b = 8'd141;  #10 
a = 8'd80; b = 8'd142;  #10 
a = 8'd80; b = 8'd143;  #10 
a = 8'd80; b = 8'd144;  #10 
a = 8'd80; b = 8'd145;  #10 
a = 8'd80; b = 8'd146;  #10 
a = 8'd80; b = 8'd147;  #10 
a = 8'd80; b = 8'd148;  #10 
a = 8'd80; b = 8'd149;  #10 
a = 8'd80; b = 8'd150;  #10 
a = 8'd80; b = 8'd151;  #10 
a = 8'd80; b = 8'd152;  #10 
a = 8'd80; b = 8'd153;  #10 
a = 8'd80; b = 8'd154;  #10 
a = 8'd80; b = 8'd155;  #10 
a = 8'd80; b = 8'd156;  #10 
a = 8'd80; b = 8'd157;  #10 
a = 8'd80; b = 8'd158;  #10 
a = 8'd80; b = 8'd159;  #10 
a = 8'd80; b = 8'd160;  #10 
a = 8'd80; b = 8'd161;  #10 
a = 8'd80; b = 8'd162;  #10 
a = 8'd80; b = 8'd163;  #10 
a = 8'd80; b = 8'd164;  #10 
a = 8'd80; b = 8'd165;  #10 
a = 8'd80; b = 8'd166;  #10 
a = 8'd80; b = 8'd167;  #10 
a = 8'd80; b = 8'd168;  #10 
a = 8'd80; b = 8'd169;  #10 
a = 8'd80; b = 8'd170;  #10 
a = 8'd80; b = 8'd171;  #10 
a = 8'd80; b = 8'd172;  #10 
a = 8'd80; b = 8'd173;  #10 
a = 8'd80; b = 8'd174;  #10 
a = 8'd80; b = 8'd175;  #10 
a = 8'd80; b = 8'd176;  #10 
a = 8'd80; b = 8'd177;  #10 
a = 8'd80; b = 8'd178;  #10 
a = 8'd80; b = 8'd179;  #10 
a = 8'd80; b = 8'd180;  #10 
a = 8'd80; b = 8'd181;  #10 
a = 8'd80; b = 8'd182;  #10 
a = 8'd80; b = 8'd183;  #10 
a = 8'd80; b = 8'd184;  #10 
a = 8'd80; b = 8'd185;  #10 
a = 8'd80; b = 8'd186;  #10 
a = 8'd80; b = 8'd187;  #10 
a = 8'd80; b = 8'd188;  #10 
a = 8'd80; b = 8'd189;  #10 
a = 8'd80; b = 8'd190;  #10 
a = 8'd80; b = 8'd191;  #10 
a = 8'd80; b = 8'd192;  #10 
a = 8'd80; b = 8'd193;  #10 
a = 8'd80; b = 8'd194;  #10 
a = 8'd80; b = 8'd195;  #10 
a = 8'd80; b = 8'd196;  #10 
a = 8'd80; b = 8'd197;  #10 
a = 8'd80; b = 8'd198;  #10 
a = 8'd80; b = 8'd199;  #10 
a = 8'd80; b = 8'd200;  #10 
a = 8'd80; b = 8'd201;  #10 
a = 8'd80; b = 8'd202;  #10 
a = 8'd80; b = 8'd203;  #10 
a = 8'd80; b = 8'd204;  #10 
a = 8'd80; b = 8'd205;  #10 
a = 8'd80; b = 8'd206;  #10 
a = 8'd80; b = 8'd207;  #10 
a = 8'd80; b = 8'd208;  #10 
a = 8'd80; b = 8'd209;  #10 
a = 8'd80; b = 8'd210;  #10 
a = 8'd80; b = 8'd211;  #10 
a = 8'd80; b = 8'd212;  #10 
a = 8'd80; b = 8'd213;  #10 
a = 8'd80; b = 8'd214;  #10 
a = 8'd80; b = 8'd215;  #10 
a = 8'd80; b = 8'd216;  #10 
a = 8'd80; b = 8'd217;  #10 
a = 8'd80; b = 8'd218;  #10 
a = 8'd80; b = 8'd219;  #10 
a = 8'd80; b = 8'd220;  #10 
a = 8'd80; b = 8'd221;  #10 
a = 8'd80; b = 8'd222;  #10 
a = 8'd80; b = 8'd223;  #10 
a = 8'd80; b = 8'd224;  #10 
a = 8'd80; b = 8'd225;  #10 
a = 8'd80; b = 8'd226;  #10 
a = 8'd80; b = 8'd227;  #10 
a = 8'd80; b = 8'd228;  #10 
a = 8'd80; b = 8'd229;  #10 
a = 8'd80; b = 8'd230;  #10 
a = 8'd80; b = 8'd231;  #10 
a = 8'd80; b = 8'd232;  #10 
a = 8'd80; b = 8'd233;  #10 
a = 8'd80; b = 8'd234;  #10 
a = 8'd80; b = 8'd235;  #10 
a = 8'd80; b = 8'd236;  #10 
a = 8'd80; b = 8'd237;  #10 
a = 8'd80; b = 8'd238;  #10 
a = 8'd80; b = 8'd239;  #10 
a = 8'd80; b = 8'd240;  #10 
a = 8'd80; b = 8'd241;  #10 
a = 8'd80; b = 8'd242;  #10 
a = 8'd80; b = 8'd243;  #10 
a = 8'd80; b = 8'd244;  #10 
a = 8'd80; b = 8'd245;  #10 
a = 8'd80; b = 8'd246;  #10 
a = 8'd80; b = 8'd247;  #10 
a = 8'd80; b = 8'd248;  #10 
a = 8'd80; b = 8'd249;  #10 
a = 8'd80; b = 8'd250;  #10 
a = 8'd80; b = 8'd251;  #10 
a = 8'd80; b = 8'd252;  #10 
a = 8'd80; b = 8'd253;  #10 
a = 8'd80; b = 8'd254;  #10 
a = 8'd80; b = 8'd255;  #10 
a = 8'd81; b = 8'd0;  #10 
a = 8'd81; b = 8'd1;  #10 
a = 8'd81; b = 8'd2;  #10 
a = 8'd81; b = 8'd3;  #10 
a = 8'd81; b = 8'd4;  #10 
a = 8'd81; b = 8'd5;  #10 
a = 8'd81; b = 8'd6;  #10 
a = 8'd81; b = 8'd7;  #10 
a = 8'd81; b = 8'd8;  #10 
a = 8'd81; b = 8'd9;  #10 
a = 8'd81; b = 8'd10;  #10 
a = 8'd81; b = 8'd11;  #10 
a = 8'd81; b = 8'd12;  #10 
a = 8'd81; b = 8'd13;  #10 
a = 8'd81; b = 8'd14;  #10 
a = 8'd81; b = 8'd15;  #10 
a = 8'd81; b = 8'd16;  #10 
a = 8'd81; b = 8'd17;  #10 
a = 8'd81; b = 8'd18;  #10 
a = 8'd81; b = 8'd19;  #10 
a = 8'd81; b = 8'd20;  #10 
a = 8'd81; b = 8'd21;  #10 
a = 8'd81; b = 8'd22;  #10 
a = 8'd81; b = 8'd23;  #10 
a = 8'd81; b = 8'd24;  #10 
a = 8'd81; b = 8'd25;  #10 
a = 8'd81; b = 8'd26;  #10 
a = 8'd81; b = 8'd27;  #10 
a = 8'd81; b = 8'd28;  #10 
a = 8'd81; b = 8'd29;  #10 
a = 8'd81; b = 8'd30;  #10 
a = 8'd81; b = 8'd31;  #10 
a = 8'd81; b = 8'd32;  #10 
a = 8'd81; b = 8'd33;  #10 
a = 8'd81; b = 8'd34;  #10 
a = 8'd81; b = 8'd35;  #10 
a = 8'd81; b = 8'd36;  #10 
a = 8'd81; b = 8'd37;  #10 
a = 8'd81; b = 8'd38;  #10 
a = 8'd81; b = 8'd39;  #10 
a = 8'd81; b = 8'd40;  #10 
a = 8'd81; b = 8'd41;  #10 
a = 8'd81; b = 8'd42;  #10 
a = 8'd81; b = 8'd43;  #10 
a = 8'd81; b = 8'd44;  #10 
a = 8'd81; b = 8'd45;  #10 
a = 8'd81; b = 8'd46;  #10 
a = 8'd81; b = 8'd47;  #10 
a = 8'd81; b = 8'd48;  #10 
a = 8'd81; b = 8'd49;  #10 
a = 8'd81; b = 8'd50;  #10 
a = 8'd81; b = 8'd51;  #10 
a = 8'd81; b = 8'd52;  #10 
a = 8'd81; b = 8'd53;  #10 
a = 8'd81; b = 8'd54;  #10 
a = 8'd81; b = 8'd55;  #10 
a = 8'd81; b = 8'd56;  #10 
a = 8'd81; b = 8'd57;  #10 
a = 8'd81; b = 8'd58;  #10 
a = 8'd81; b = 8'd59;  #10 
a = 8'd81; b = 8'd60;  #10 
a = 8'd81; b = 8'd61;  #10 
a = 8'd81; b = 8'd62;  #10 
a = 8'd81; b = 8'd63;  #10 
a = 8'd81; b = 8'd64;  #10 
a = 8'd81; b = 8'd65;  #10 
a = 8'd81; b = 8'd66;  #10 
a = 8'd81; b = 8'd67;  #10 
a = 8'd81; b = 8'd68;  #10 
a = 8'd81; b = 8'd69;  #10 
a = 8'd81; b = 8'd70;  #10 
a = 8'd81; b = 8'd71;  #10 
a = 8'd81; b = 8'd72;  #10 
a = 8'd81; b = 8'd73;  #10 
a = 8'd81; b = 8'd74;  #10 
a = 8'd81; b = 8'd75;  #10 
a = 8'd81; b = 8'd76;  #10 
a = 8'd81; b = 8'd77;  #10 
a = 8'd81; b = 8'd78;  #10 
a = 8'd81; b = 8'd79;  #10 
a = 8'd81; b = 8'd80;  #10 
a = 8'd81; b = 8'd81;  #10 
a = 8'd81; b = 8'd82;  #10 
a = 8'd81; b = 8'd83;  #10 
a = 8'd81; b = 8'd84;  #10 
a = 8'd81; b = 8'd85;  #10 
a = 8'd81; b = 8'd86;  #10 
a = 8'd81; b = 8'd87;  #10 
a = 8'd81; b = 8'd88;  #10 
a = 8'd81; b = 8'd89;  #10 
a = 8'd81; b = 8'd90;  #10 
a = 8'd81; b = 8'd91;  #10 
a = 8'd81; b = 8'd92;  #10 
a = 8'd81; b = 8'd93;  #10 
a = 8'd81; b = 8'd94;  #10 
a = 8'd81; b = 8'd95;  #10 
a = 8'd81; b = 8'd96;  #10 
a = 8'd81; b = 8'd97;  #10 
a = 8'd81; b = 8'd98;  #10 
a = 8'd81; b = 8'd99;  #10 
a = 8'd81; b = 8'd100;  #10 
a = 8'd81; b = 8'd101;  #10 
a = 8'd81; b = 8'd102;  #10 
a = 8'd81; b = 8'd103;  #10 
a = 8'd81; b = 8'd104;  #10 
a = 8'd81; b = 8'd105;  #10 
a = 8'd81; b = 8'd106;  #10 
a = 8'd81; b = 8'd107;  #10 
a = 8'd81; b = 8'd108;  #10 
a = 8'd81; b = 8'd109;  #10 
a = 8'd81; b = 8'd110;  #10 
a = 8'd81; b = 8'd111;  #10 
a = 8'd81; b = 8'd112;  #10 
a = 8'd81; b = 8'd113;  #10 
a = 8'd81; b = 8'd114;  #10 
a = 8'd81; b = 8'd115;  #10 
a = 8'd81; b = 8'd116;  #10 
a = 8'd81; b = 8'd117;  #10 
a = 8'd81; b = 8'd118;  #10 
a = 8'd81; b = 8'd119;  #10 
a = 8'd81; b = 8'd120;  #10 
a = 8'd81; b = 8'd121;  #10 
a = 8'd81; b = 8'd122;  #10 
a = 8'd81; b = 8'd123;  #10 
a = 8'd81; b = 8'd124;  #10 
a = 8'd81; b = 8'd125;  #10 
a = 8'd81; b = 8'd126;  #10 
a = 8'd81; b = 8'd127;  #10 
a = 8'd81; b = 8'd128;  #10 
a = 8'd81; b = 8'd129;  #10 
a = 8'd81; b = 8'd130;  #10 
a = 8'd81; b = 8'd131;  #10 
a = 8'd81; b = 8'd132;  #10 
a = 8'd81; b = 8'd133;  #10 
a = 8'd81; b = 8'd134;  #10 
a = 8'd81; b = 8'd135;  #10 
a = 8'd81; b = 8'd136;  #10 
a = 8'd81; b = 8'd137;  #10 
a = 8'd81; b = 8'd138;  #10 
a = 8'd81; b = 8'd139;  #10 
a = 8'd81; b = 8'd140;  #10 
a = 8'd81; b = 8'd141;  #10 
a = 8'd81; b = 8'd142;  #10 
a = 8'd81; b = 8'd143;  #10 
a = 8'd81; b = 8'd144;  #10 
a = 8'd81; b = 8'd145;  #10 
a = 8'd81; b = 8'd146;  #10 
a = 8'd81; b = 8'd147;  #10 
a = 8'd81; b = 8'd148;  #10 
a = 8'd81; b = 8'd149;  #10 
a = 8'd81; b = 8'd150;  #10 
a = 8'd81; b = 8'd151;  #10 
a = 8'd81; b = 8'd152;  #10 
a = 8'd81; b = 8'd153;  #10 
a = 8'd81; b = 8'd154;  #10 
a = 8'd81; b = 8'd155;  #10 
a = 8'd81; b = 8'd156;  #10 
a = 8'd81; b = 8'd157;  #10 
a = 8'd81; b = 8'd158;  #10 
a = 8'd81; b = 8'd159;  #10 
a = 8'd81; b = 8'd160;  #10 
a = 8'd81; b = 8'd161;  #10 
a = 8'd81; b = 8'd162;  #10 
a = 8'd81; b = 8'd163;  #10 
a = 8'd81; b = 8'd164;  #10 
a = 8'd81; b = 8'd165;  #10 
a = 8'd81; b = 8'd166;  #10 
a = 8'd81; b = 8'd167;  #10 
a = 8'd81; b = 8'd168;  #10 
a = 8'd81; b = 8'd169;  #10 
a = 8'd81; b = 8'd170;  #10 
a = 8'd81; b = 8'd171;  #10 
a = 8'd81; b = 8'd172;  #10 
a = 8'd81; b = 8'd173;  #10 
a = 8'd81; b = 8'd174;  #10 
a = 8'd81; b = 8'd175;  #10 
a = 8'd81; b = 8'd176;  #10 
a = 8'd81; b = 8'd177;  #10 
a = 8'd81; b = 8'd178;  #10 
a = 8'd81; b = 8'd179;  #10 
a = 8'd81; b = 8'd180;  #10 
a = 8'd81; b = 8'd181;  #10 
a = 8'd81; b = 8'd182;  #10 
a = 8'd81; b = 8'd183;  #10 
a = 8'd81; b = 8'd184;  #10 
a = 8'd81; b = 8'd185;  #10 
a = 8'd81; b = 8'd186;  #10 
a = 8'd81; b = 8'd187;  #10 
a = 8'd81; b = 8'd188;  #10 
a = 8'd81; b = 8'd189;  #10 
a = 8'd81; b = 8'd190;  #10 
a = 8'd81; b = 8'd191;  #10 
a = 8'd81; b = 8'd192;  #10 
a = 8'd81; b = 8'd193;  #10 
a = 8'd81; b = 8'd194;  #10 
a = 8'd81; b = 8'd195;  #10 
a = 8'd81; b = 8'd196;  #10 
a = 8'd81; b = 8'd197;  #10 
a = 8'd81; b = 8'd198;  #10 
a = 8'd81; b = 8'd199;  #10 
a = 8'd81; b = 8'd200;  #10 
a = 8'd81; b = 8'd201;  #10 
a = 8'd81; b = 8'd202;  #10 
a = 8'd81; b = 8'd203;  #10 
a = 8'd81; b = 8'd204;  #10 
a = 8'd81; b = 8'd205;  #10 
a = 8'd81; b = 8'd206;  #10 
a = 8'd81; b = 8'd207;  #10 
a = 8'd81; b = 8'd208;  #10 
a = 8'd81; b = 8'd209;  #10 
a = 8'd81; b = 8'd210;  #10 
a = 8'd81; b = 8'd211;  #10 
a = 8'd81; b = 8'd212;  #10 
a = 8'd81; b = 8'd213;  #10 
a = 8'd81; b = 8'd214;  #10 
a = 8'd81; b = 8'd215;  #10 
a = 8'd81; b = 8'd216;  #10 
a = 8'd81; b = 8'd217;  #10 
a = 8'd81; b = 8'd218;  #10 
a = 8'd81; b = 8'd219;  #10 
a = 8'd81; b = 8'd220;  #10 
a = 8'd81; b = 8'd221;  #10 
a = 8'd81; b = 8'd222;  #10 
a = 8'd81; b = 8'd223;  #10 
a = 8'd81; b = 8'd224;  #10 
a = 8'd81; b = 8'd225;  #10 
a = 8'd81; b = 8'd226;  #10 
a = 8'd81; b = 8'd227;  #10 
a = 8'd81; b = 8'd228;  #10 
a = 8'd81; b = 8'd229;  #10 
a = 8'd81; b = 8'd230;  #10 
a = 8'd81; b = 8'd231;  #10 
a = 8'd81; b = 8'd232;  #10 
a = 8'd81; b = 8'd233;  #10 
a = 8'd81; b = 8'd234;  #10 
a = 8'd81; b = 8'd235;  #10 
a = 8'd81; b = 8'd236;  #10 
a = 8'd81; b = 8'd237;  #10 
a = 8'd81; b = 8'd238;  #10 
a = 8'd81; b = 8'd239;  #10 
a = 8'd81; b = 8'd240;  #10 
a = 8'd81; b = 8'd241;  #10 
a = 8'd81; b = 8'd242;  #10 
a = 8'd81; b = 8'd243;  #10 
a = 8'd81; b = 8'd244;  #10 
a = 8'd81; b = 8'd245;  #10 
a = 8'd81; b = 8'd246;  #10 
a = 8'd81; b = 8'd247;  #10 
a = 8'd81; b = 8'd248;  #10 
a = 8'd81; b = 8'd249;  #10 
a = 8'd81; b = 8'd250;  #10 
a = 8'd81; b = 8'd251;  #10 
a = 8'd81; b = 8'd252;  #10 
a = 8'd81; b = 8'd253;  #10 
a = 8'd81; b = 8'd254;  #10 
a = 8'd81; b = 8'd255;  #10 
a = 8'd82; b = 8'd0;  #10 
a = 8'd82; b = 8'd1;  #10 
a = 8'd82; b = 8'd2;  #10 
a = 8'd82; b = 8'd3;  #10 
a = 8'd82; b = 8'd4;  #10 
a = 8'd82; b = 8'd5;  #10 
a = 8'd82; b = 8'd6;  #10 
a = 8'd82; b = 8'd7;  #10 
a = 8'd82; b = 8'd8;  #10 
a = 8'd82; b = 8'd9;  #10 
a = 8'd82; b = 8'd10;  #10 
a = 8'd82; b = 8'd11;  #10 
a = 8'd82; b = 8'd12;  #10 
a = 8'd82; b = 8'd13;  #10 
a = 8'd82; b = 8'd14;  #10 
a = 8'd82; b = 8'd15;  #10 
a = 8'd82; b = 8'd16;  #10 
a = 8'd82; b = 8'd17;  #10 
a = 8'd82; b = 8'd18;  #10 
a = 8'd82; b = 8'd19;  #10 
a = 8'd82; b = 8'd20;  #10 
a = 8'd82; b = 8'd21;  #10 
a = 8'd82; b = 8'd22;  #10 
a = 8'd82; b = 8'd23;  #10 
a = 8'd82; b = 8'd24;  #10 
a = 8'd82; b = 8'd25;  #10 
a = 8'd82; b = 8'd26;  #10 
a = 8'd82; b = 8'd27;  #10 
a = 8'd82; b = 8'd28;  #10 
a = 8'd82; b = 8'd29;  #10 
a = 8'd82; b = 8'd30;  #10 
a = 8'd82; b = 8'd31;  #10 
a = 8'd82; b = 8'd32;  #10 
a = 8'd82; b = 8'd33;  #10 
a = 8'd82; b = 8'd34;  #10 
a = 8'd82; b = 8'd35;  #10 
a = 8'd82; b = 8'd36;  #10 
a = 8'd82; b = 8'd37;  #10 
a = 8'd82; b = 8'd38;  #10 
a = 8'd82; b = 8'd39;  #10 
a = 8'd82; b = 8'd40;  #10 
a = 8'd82; b = 8'd41;  #10 
a = 8'd82; b = 8'd42;  #10 
a = 8'd82; b = 8'd43;  #10 
a = 8'd82; b = 8'd44;  #10 
a = 8'd82; b = 8'd45;  #10 
a = 8'd82; b = 8'd46;  #10 
a = 8'd82; b = 8'd47;  #10 
a = 8'd82; b = 8'd48;  #10 
a = 8'd82; b = 8'd49;  #10 
a = 8'd82; b = 8'd50;  #10 
a = 8'd82; b = 8'd51;  #10 
a = 8'd82; b = 8'd52;  #10 
a = 8'd82; b = 8'd53;  #10 
a = 8'd82; b = 8'd54;  #10 
a = 8'd82; b = 8'd55;  #10 
a = 8'd82; b = 8'd56;  #10 
a = 8'd82; b = 8'd57;  #10 
a = 8'd82; b = 8'd58;  #10 
a = 8'd82; b = 8'd59;  #10 
a = 8'd82; b = 8'd60;  #10 
a = 8'd82; b = 8'd61;  #10 
a = 8'd82; b = 8'd62;  #10 
a = 8'd82; b = 8'd63;  #10 
a = 8'd82; b = 8'd64;  #10 
a = 8'd82; b = 8'd65;  #10 
a = 8'd82; b = 8'd66;  #10 
a = 8'd82; b = 8'd67;  #10 
a = 8'd82; b = 8'd68;  #10 
a = 8'd82; b = 8'd69;  #10 
a = 8'd82; b = 8'd70;  #10 
a = 8'd82; b = 8'd71;  #10 
a = 8'd82; b = 8'd72;  #10 
a = 8'd82; b = 8'd73;  #10 
a = 8'd82; b = 8'd74;  #10 
a = 8'd82; b = 8'd75;  #10 
a = 8'd82; b = 8'd76;  #10 
a = 8'd82; b = 8'd77;  #10 
a = 8'd82; b = 8'd78;  #10 
a = 8'd82; b = 8'd79;  #10 
a = 8'd82; b = 8'd80;  #10 
a = 8'd82; b = 8'd81;  #10 
a = 8'd82; b = 8'd82;  #10 
a = 8'd82; b = 8'd83;  #10 
a = 8'd82; b = 8'd84;  #10 
a = 8'd82; b = 8'd85;  #10 
a = 8'd82; b = 8'd86;  #10 
a = 8'd82; b = 8'd87;  #10 
a = 8'd82; b = 8'd88;  #10 
a = 8'd82; b = 8'd89;  #10 
a = 8'd82; b = 8'd90;  #10 
a = 8'd82; b = 8'd91;  #10 
a = 8'd82; b = 8'd92;  #10 
a = 8'd82; b = 8'd93;  #10 
a = 8'd82; b = 8'd94;  #10 
a = 8'd82; b = 8'd95;  #10 
a = 8'd82; b = 8'd96;  #10 
a = 8'd82; b = 8'd97;  #10 
a = 8'd82; b = 8'd98;  #10 
a = 8'd82; b = 8'd99;  #10 
a = 8'd82; b = 8'd100;  #10 
a = 8'd82; b = 8'd101;  #10 
a = 8'd82; b = 8'd102;  #10 
a = 8'd82; b = 8'd103;  #10 
a = 8'd82; b = 8'd104;  #10 
a = 8'd82; b = 8'd105;  #10 
a = 8'd82; b = 8'd106;  #10 
a = 8'd82; b = 8'd107;  #10 
a = 8'd82; b = 8'd108;  #10 
a = 8'd82; b = 8'd109;  #10 
a = 8'd82; b = 8'd110;  #10 
a = 8'd82; b = 8'd111;  #10 
a = 8'd82; b = 8'd112;  #10 
a = 8'd82; b = 8'd113;  #10 
a = 8'd82; b = 8'd114;  #10 
a = 8'd82; b = 8'd115;  #10 
a = 8'd82; b = 8'd116;  #10 
a = 8'd82; b = 8'd117;  #10 
a = 8'd82; b = 8'd118;  #10 
a = 8'd82; b = 8'd119;  #10 
a = 8'd82; b = 8'd120;  #10 
a = 8'd82; b = 8'd121;  #10 
a = 8'd82; b = 8'd122;  #10 
a = 8'd82; b = 8'd123;  #10 
a = 8'd82; b = 8'd124;  #10 
a = 8'd82; b = 8'd125;  #10 
a = 8'd82; b = 8'd126;  #10 
a = 8'd82; b = 8'd127;  #10 
a = 8'd82; b = 8'd128;  #10 
a = 8'd82; b = 8'd129;  #10 
a = 8'd82; b = 8'd130;  #10 
a = 8'd82; b = 8'd131;  #10 
a = 8'd82; b = 8'd132;  #10 
a = 8'd82; b = 8'd133;  #10 
a = 8'd82; b = 8'd134;  #10 
a = 8'd82; b = 8'd135;  #10 
a = 8'd82; b = 8'd136;  #10 
a = 8'd82; b = 8'd137;  #10 
a = 8'd82; b = 8'd138;  #10 
a = 8'd82; b = 8'd139;  #10 
a = 8'd82; b = 8'd140;  #10 
a = 8'd82; b = 8'd141;  #10 
a = 8'd82; b = 8'd142;  #10 
a = 8'd82; b = 8'd143;  #10 
a = 8'd82; b = 8'd144;  #10 
a = 8'd82; b = 8'd145;  #10 
a = 8'd82; b = 8'd146;  #10 
a = 8'd82; b = 8'd147;  #10 
a = 8'd82; b = 8'd148;  #10 
a = 8'd82; b = 8'd149;  #10 
a = 8'd82; b = 8'd150;  #10 
a = 8'd82; b = 8'd151;  #10 
a = 8'd82; b = 8'd152;  #10 
a = 8'd82; b = 8'd153;  #10 
a = 8'd82; b = 8'd154;  #10 
a = 8'd82; b = 8'd155;  #10 
a = 8'd82; b = 8'd156;  #10 
a = 8'd82; b = 8'd157;  #10 
a = 8'd82; b = 8'd158;  #10 
a = 8'd82; b = 8'd159;  #10 
a = 8'd82; b = 8'd160;  #10 
a = 8'd82; b = 8'd161;  #10 
a = 8'd82; b = 8'd162;  #10 
a = 8'd82; b = 8'd163;  #10 
a = 8'd82; b = 8'd164;  #10 
a = 8'd82; b = 8'd165;  #10 
a = 8'd82; b = 8'd166;  #10 
a = 8'd82; b = 8'd167;  #10 
a = 8'd82; b = 8'd168;  #10 
a = 8'd82; b = 8'd169;  #10 
a = 8'd82; b = 8'd170;  #10 
a = 8'd82; b = 8'd171;  #10 
a = 8'd82; b = 8'd172;  #10 
a = 8'd82; b = 8'd173;  #10 
a = 8'd82; b = 8'd174;  #10 
a = 8'd82; b = 8'd175;  #10 
a = 8'd82; b = 8'd176;  #10 
a = 8'd82; b = 8'd177;  #10 
a = 8'd82; b = 8'd178;  #10 
a = 8'd82; b = 8'd179;  #10 
a = 8'd82; b = 8'd180;  #10 
a = 8'd82; b = 8'd181;  #10 
a = 8'd82; b = 8'd182;  #10 
a = 8'd82; b = 8'd183;  #10 
a = 8'd82; b = 8'd184;  #10 
a = 8'd82; b = 8'd185;  #10 
a = 8'd82; b = 8'd186;  #10 
a = 8'd82; b = 8'd187;  #10 
a = 8'd82; b = 8'd188;  #10 
a = 8'd82; b = 8'd189;  #10 
a = 8'd82; b = 8'd190;  #10 
a = 8'd82; b = 8'd191;  #10 
a = 8'd82; b = 8'd192;  #10 
a = 8'd82; b = 8'd193;  #10 
a = 8'd82; b = 8'd194;  #10 
a = 8'd82; b = 8'd195;  #10 
a = 8'd82; b = 8'd196;  #10 
a = 8'd82; b = 8'd197;  #10 
a = 8'd82; b = 8'd198;  #10 
a = 8'd82; b = 8'd199;  #10 
a = 8'd82; b = 8'd200;  #10 
a = 8'd82; b = 8'd201;  #10 
a = 8'd82; b = 8'd202;  #10 
a = 8'd82; b = 8'd203;  #10 
a = 8'd82; b = 8'd204;  #10 
a = 8'd82; b = 8'd205;  #10 
a = 8'd82; b = 8'd206;  #10 
a = 8'd82; b = 8'd207;  #10 
a = 8'd82; b = 8'd208;  #10 
a = 8'd82; b = 8'd209;  #10 
a = 8'd82; b = 8'd210;  #10 
a = 8'd82; b = 8'd211;  #10 
a = 8'd82; b = 8'd212;  #10 
a = 8'd82; b = 8'd213;  #10 
a = 8'd82; b = 8'd214;  #10 
a = 8'd82; b = 8'd215;  #10 
a = 8'd82; b = 8'd216;  #10 
a = 8'd82; b = 8'd217;  #10 
a = 8'd82; b = 8'd218;  #10 
a = 8'd82; b = 8'd219;  #10 
a = 8'd82; b = 8'd220;  #10 
a = 8'd82; b = 8'd221;  #10 
a = 8'd82; b = 8'd222;  #10 
a = 8'd82; b = 8'd223;  #10 
a = 8'd82; b = 8'd224;  #10 
a = 8'd82; b = 8'd225;  #10 
a = 8'd82; b = 8'd226;  #10 
a = 8'd82; b = 8'd227;  #10 
a = 8'd82; b = 8'd228;  #10 
a = 8'd82; b = 8'd229;  #10 
a = 8'd82; b = 8'd230;  #10 
a = 8'd82; b = 8'd231;  #10 
a = 8'd82; b = 8'd232;  #10 
a = 8'd82; b = 8'd233;  #10 
a = 8'd82; b = 8'd234;  #10 
a = 8'd82; b = 8'd235;  #10 
a = 8'd82; b = 8'd236;  #10 
a = 8'd82; b = 8'd237;  #10 
a = 8'd82; b = 8'd238;  #10 
a = 8'd82; b = 8'd239;  #10 
a = 8'd82; b = 8'd240;  #10 
a = 8'd82; b = 8'd241;  #10 
a = 8'd82; b = 8'd242;  #10 
a = 8'd82; b = 8'd243;  #10 
a = 8'd82; b = 8'd244;  #10 
a = 8'd82; b = 8'd245;  #10 
a = 8'd82; b = 8'd246;  #10 
a = 8'd82; b = 8'd247;  #10 
a = 8'd82; b = 8'd248;  #10 
a = 8'd82; b = 8'd249;  #10 
a = 8'd82; b = 8'd250;  #10 
a = 8'd82; b = 8'd251;  #10 
a = 8'd82; b = 8'd252;  #10 
a = 8'd82; b = 8'd253;  #10 
a = 8'd82; b = 8'd254;  #10 
a = 8'd82; b = 8'd255;  #10 
a = 8'd83; b = 8'd0;  #10 
a = 8'd83; b = 8'd1;  #10 
a = 8'd83; b = 8'd2;  #10 
a = 8'd83; b = 8'd3;  #10 
a = 8'd83; b = 8'd4;  #10 
a = 8'd83; b = 8'd5;  #10 
a = 8'd83; b = 8'd6;  #10 
a = 8'd83; b = 8'd7;  #10 
a = 8'd83; b = 8'd8;  #10 
a = 8'd83; b = 8'd9;  #10 
a = 8'd83; b = 8'd10;  #10 
a = 8'd83; b = 8'd11;  #10 
a = 8'd83; b = 8'd12;  #10 
a = 8'd83; b = 8'd13;  #10 
a = 8'd83; b = 8'd14;  #10 
a = 8'd83; b = 8'd15;  #10 
a = 8'd83; b = 8'd16;  #10 
a = 8'd83; b = 8'd17;  #10 
a = 8'd83; b = 8'd18;  #10 
a = 8'd83; b = 8'd19;  #10 
a = 8'd83; b = 8'd20;  #10 
a = 8'd83; b = 8'd21;  #10 
a = 8'd83; b = 8'd22;  #10 
a = 8'd83; b = 8'd23;  #10 
a = 8'd83; b = 8'd24;  #10 
a = 8'd83; b = 8'd25;  #10 
a = 8'd83; b = 8'd26;  #10 
a = 8'd83; b = 8'd27;  #10 
a = 8'd83; b = 8'd28;  #10 
a = 8'd83; b = 8'd29;  #10 
a = 8'd83; b = 8'd30;  #10 
a = 8'd83; b = 8'd31;  #10 
a = 8'd83; b = 8'd32;  #10 
a = 8'd83; b = 8'd33;  #10 
a = 8'd83; b = 8'd34;  #10 
a = 8'd83; b = 8'd35;  #10 
a = 8'd83; b = 8'd36;  #10 
a = 8'd83; b = 8'd37;  #10 
a = 8'd83; b = 8'd38;  #10 
a = 8'd83; b = 8'd39;  #10 
a = 8'd83; b = 8'd40;  #10 
a = 8'd83; b = 8'd41;  #10 
a = 8'd83; b = 8'd42;  #10 
a = 8'd83; b = 8'd43;  #10 
a = 8'd83; b = 8'd44;  #10 
a = 8'd83; b = 8'd45;  #10 
a = 8'd83; b = 8'd46;  #10 
a = 8'd83; b = 8'd47;  #10 
a = 8'd83; b = 8'd48;  #10 
a = 8'd83; b = 8'd49;  #10 
a = 8'd83; b = 8'd50;  #10 
a = 8'd83; b = 8'd51;  #10 
a = 8'd83; b = 8'd52;  #10 
a = 8'd83; b = 8'd53;  #10 
a = 8'd83; b = 8'd54;  #10 
a = 8'd83; b = 8'd55;  #10 
a = 8'd83; b = 8'd56;  #10 
a = 8'd83; b = 8'd57;  #10 
a = 8'd83; b = 8'd58;  #10 
a = 8'd83; b = 8'd59;  #10 
a = 8'd83; b = 8'd60;  #10 
a = 8'd83; b = 8'd61;  #10 
a = 8'd83; b = 8'd62;  #10 
a = 8'd83; b = 8'd63;  #10 
a = 8'd83; b = 8'd64;  #10 
a = 8'd83; b = 8'd65;  #10 
a = 8'd83; b = 8'd66;  #10 
a = 8'd83; b = 8'd67;  #10 
a = 8'd83; b = 8'd68;  #10 
a = 8'd83; b = 8'd69;  #10 
a = 8'd83; b = 8'd70;  #10 
a = 8'd83; b = 8'd71;  #10 
a = 8'd83; b = 8'd72;  #10 
a = 8'd83; b = 8'd73;  #10 
a = 8'd83; b = 8'd74;  #10 
a = 8'd83; b = 8'd75;  #10 
a = 8'd83; b = 8'd76;  #10 
a = 8'd83; b = 8'd77;  #10 
a = 8'd83; b = 8'd78;  #10 
a = 8'd83; b = 8'd79;  #10 
a = 8'd83; b = 8'd80;  #10 
a = 8'd83; b = 8'd81;  #10 
a = 8'd83; b = 8'd82;  #10 
a = 8'd83; b = 8'd83;  #10 
a = 8'd83; b = 8'd84;  #10 
a = 8'd83; b = 8'd85;  #10 
a = 8'd83; b = 8'd86;  #10 
a = 8'd83; b = 8'd87;  #10 
a = 8'd83; b = 8'd88;  #10 
a = 8'd83; b = 8'd89;  #10 
a = 8'd83; b = 8'd90;  #10 
a = 8'd83; b = 8'd91;  #10 
a = 8'd83; b = 8'd92;  #10 
a = 8'd83; b = 8'd93;  #10 
a = 8'd83; b = 8'd94;  #10 
a = 8'd83; b = 8'd95;  #10 
a = 8'd83; b = 8'd96;  #10 
a = 8'd83; b = 8'd97;  #10 
a = 8'd83; b = 8'd98;  #10 
a = 8'd83; b = 8'd99;  #10 
a = 8'd83; b = 8'd100;  #10 
a = 8'd83; b = 8'd101;  #10 
a = 8'd83; b = 8'd102;  #10 
a = 8'd83; b = 8'd103;  #10 
a = 8'd83; b = 8'd104;  #10 
a = 8'd83; b = 8'd105;  #10 
a = 8'd83; b = 8'd106;  #10 
a = 8'd83; b = 8'd107;  #10 
a = 8'd83; b = 8'd108;  #10 
a = 8'd83; b = 8'd109;  #10 
a = 8'd83; b = 8'd110;  #10 
a = 8'd83; b = 8'd111;  #10 
a = 8'd83; b = 8'd112;  #10 
a = 8'd83; b = 8'd113;  #10 
a = 8'd83; b = 8'd114;  #10 
a = 8'd83; b = 8'd115;  #10 
a = 8'd83; b = 8'd116;  #10 
a = 8'd83; b = 8'd117;  #10 
a = 8'd83; b = 8'd118;  #10 
a = 8'd83; b = 8'd119;  #10 
a = 8'd83; b = 8'd120;  #10 
a = 8'd83; b = 8'd121;  #10 
a = 8'd83; b = 8'd122;  #10 
a = 8'd83; b = 8'd123;  #10 
a = 8'd83; b = 8'd124;  #10 
a = 8'd83; b = 8'd125;  #10 
a = 8'd83; b = 8'd126;  #10 
a = 8'd83; b = 8'd127;  #10 
a = 8'd83; b = 8'd128;  #10 
a = 8'd83; b = 8'd129;  #10 
a = 8'd83; b = 8'd130;  #10 
a = 8'd83; b = 8'd131;  #10 
a = 8'd83; b = 8'd132;  #10 
a = 8'd83; b = 8'd133;  #10 
a = 8'd83; b = 8'd134;  #10 
a = 8'd83; b = 8'd135;  #10 
a = 8'd83; b = 8'd136;  #10 
a = 8'd83; b = 8'd137;  #10 
a = 8'd83; b = 8'd138;  #10 
a = 8'd83; b = 8'd139;  #10 
a = 8'd83; b = 8'd140;  #10 
a = 8'd83; b = 8'd141;  #10 
a = 8'd83; b = 8'd142;  #10 
a = 8'd83; b = 8'd143;  #10 
a = 8'd83; b = 8'd144;  #10 
a = 8'd83; b = 8'd145;  #10 
a = 8'd83; b = 8'd146;  #10 
a = 8'd83; b = 8'd147;  #10 
a = 8'd83; b = 8'd148;  #10 
a = 8'd83; b = 8'd149;  #10 
a = 8'd83; b = 8'd150;  #10 
a = 8'd83; b = 8'd151;  #10 
a = 8'd83; b = 8'd152;  #10 
a = 8'd83; b = 8'd153;  #10 
a = 8'd83; b = 8'd154;  #10 
a = 8'd83; b = 8'd155;  #10 
a = 8'd83; b = 8'd156;  #10 
a = 8'd83; b = 8'd157;  #10 
a = 8'd83; b = 8'd158;  #10 
a = 8'd83; b = 8'd159;  #10 
a = 8'd83; b = 8'd160;  #10 
a = 8'd83; b = 8'd161;  #10 
a = 8'd83; b = 8'd162;  #10 
a = 8'd83; b = 8'd163;  #10 
a = 8'd83; b = 8'd164;  #10 
a = 8'd83; b = 8'd165;  #10 
a = 8'd83; b = 8'd166;  #10 
a = 8'd83; b = 8'd167;  #10 
a = 8'd83; b = 8'd168;  #10 
a = 8'd83; b = 8'd169;  #10 
a = 8'd83; b = 8'd170;  #10 
a = 8'd83; b = 8'd171;  #10 
a = 8'd83; b = 8'd172;  #10 
a = 8'd83; b = 8'd173;  #10 
a = 8'd83; b = 8'd174;  #10 
a = 8'd83; b = 8'd175;  #10 
a = 8'd83; b = 8'd176;  #10 
a = 8'd83; b = 8'd177;  #10 
a = 8'd83; b = 8'd178;  #10 
a = 8'd83; b = 8'd179;  #10 
a = 8'd83; b = 8'd180;  #10 
a = 8'd83; b = 8'd181;  #10 
a = 8'd83; b = 8'd182;  #10 
a = 8'd83; b = 8'd183;  #10 
a = 8'd83; b = 8'd184;  #10 
a = 8'd83; b = 8'd185;  #10 
a = 8'd83; b = 8'd186;  #10 
a = 8'd83; b = 8'd187;  #10 
a = 8'd83; b = 8'd188;  #10 
a = 8'd83; b = 8'd189;  #10 
a = 8'd83; b = 8'd190;  #10 
a = 8'd83; b = 8'd191;  #10 
a = 8'd83; b = 8'd192;  #10 
a = 8'd83; b = 8'd193;  #10 
a = 8'd83; b = 8'd194;  #10 
a = 8'd83; b = 8'd195;  #10 
a = 8'd83; b = 8'd196;  #10 
a = 8'd83; b = 8'd197;  #10 
a = 8'd83; b = 8'd198;  #10 
a = 8'd83; b = 8'd199;  #10 
a = 8'd83; b = 8'd200;  #10 
a = 8'd83; b = 8'd201;  #10 
a = 8'd83; b = 8'd202;  #10 
a = 8'd83; b = 8'd203;  #10 
a = 8'd83; b = 8'd204;  #10 
a = 8'd83; b = 8'd205;  #10 
a = 8'd83; b = 8'd206;  #10 
a = 8'd83; b = 8'd207;  #10 
a = 8'd83; b = 8'd208;  #10 
a = 8'd83; b = 8'd209;  #10 
a = 8'd83; b = 8'd210;  #10 
a = 8'd83; b = 8'd211;  #10 
a = 8'd83; b = 8'd212;  #10 
a = 8'd83; b = 8'd213;  #10 
a = 8'd83; b = 8'd214;  #10 
a = 8'd83; b = 8'd215;  #10 
a = 8'd83; b = 8'd216;  #10 
a = 8'd83; b = 8'd217;  #10 
a = 8'd83; b = 8'd218;  #10 
a = 8'd83; b = 8'd219;  #10 
a = 8'd83; b = 8'd220;  #10 
a = 8'd83; b = 8'd221;  #10 
a = 8'd83; b = 8'd222;  #10 
a = 8'd83; b = 8'd223;  #10 
a = 8'd83; b = 8'd224;  #10 
a = 8'd83; b = 8'd225;  #10 
a = 8'd83; b = 8'd226;  #10 
a = 8'd83; b = 8'd227;  #10 
a = 8'd83; b = 8'd228;  #10 
a = 8'd83; b = 8'd229;  #10 
a = 8'd83; b = 8'd230;  #10 
a = 8'd83; b = 8'd231;  #10 
a = 8'd83; b = 8'd232;  #10 
a = 8'd83; b = 8'd233;  #10 
a = 8'd83; b = 8'd234;  #10 
a = 8'd83; b = 8'd235;  #10 
a = 8'd83; b = 8'd236;  #10 
a = 8'd83; b = 8'd237;  #10 
a = 8'd83; b = 8'd238;  #10 
a = 8'd83; b = 8'd239;  #10 
a = 8'd83; b = 8'd240;  #10 
a = 8'd83; b = 8'd241;  #10 
a = 8'd83; b = 8'd242;  #10 
a = 8'd83; b = 8'd243;  #10 
a = 8'd83; b = 8'd244;  #10 
a = 8'd83; b = 8'd245;  #10 
a = 8'd83; b = 8'd246;  #10 
a = 8'd83; b = 8'd247;  #10 
a = 8'd83; b = 8'd248;  #10 
a = 8'd83; b = 8'd249;  #10 
a = 8'd83; b = 8'd250;  #10 
a = 8'd83; b = 8'd251;  #10 
a = 8'd83; b = 8'd252;  #10 
a = 8'd83; b = 8'd253;  #10 
a = 8'd83; b = 8'd254;  #10 
a = 8'd83; b = 8'd255;  #10 
a = 8'd84; b = 8'd0;  #10 
a = 8'd84; b = 8'd1;  #10 
a = 8'd84; b = 8'd2;  #10 
a = 8'd84; b = 8'd3;  #10 
a = 8'd84; b = 8'd4;  #10 
a = 8'd84; b = 8'd5;  #10 
a = 8'd84; b = 8'd6;  #10 
a = 8'd84; b = 8'd7;  #10 
a = 8'd84; b = 8'd8;  #10 
a = 8'd84; b = 8'd9;  #10 
a = 8'd84; b = 8'd10;  #10 
a = 8'd84; b = 8'd11;  #10 
a = 8'd84; b = 8'd12;  #10 
a = 8'd84; b = 8'd13;  #10 
a = 8'd84; b = 8'd14;  #10 
a = 8'd84; b = 8'd15;  #10 
a = 8'd84; b = 8'd16;  #10 
a = 8'd84; b = 8'd17;  #10 
a = 8'd84; b = 8'd18;  #10 
a = 8'd84; b = 8'd19;  #10 
a = 8'd84; b = 8'd20;  #10 
a = 8'd84; b = 8'd21;  #10 
a = 8'd84; b = 8'd22;  #10 
a = 8'd84; b = 8'd23;  #10 
a = 8'd84; b = 8'd24;  #10 
a = 8'd84; b = 8'd25;  #10 
a = 8'd84; b = 8'd26;  #10 
a = 8'd84; b = 8'd27;  #10 
a = 8'd84; b = 8'd28;  #10 
a = 8'd84; b = 8'd29;  #10 
a = 8'd84; b = 8'd30;  #10 
a = 8'd84; b = 8'd31;  #10 
a = 8'd84; b = 8'd32;  #10 
a = 8'd84; b = 8'd33;  #10 
a = 8'd84; b = 8'd34;  #10 
a = 8'd84; b = 8'd35;  #10 
a = 8'd84; b = 8'd36;  #10 
a = 8'd84; b = 8'd37;  #10 
a = 8'd84; b = 8'd38;  #10 
a = 8'd84; b = 8'd39;  #10 
a = 8'd84; b = 8'd40;  #10 
a = 8'd84; b = 8'd41;  #10 
a = 8'd84; b = 8'd42;  #10 
a = 8'd84; b = 8'd43;  #10 
a = 8'd84; b = 8'd44;  #10 
a = 8'd84; b = 8'd45;  #10 
a = 8'd84; b = 8'd46;  #10 
a = 8'd84; b = 8'd47;  #10 
a = 8'd84; b = 8'd48;  #10 
a = 8'd84; b = 8'd49;  #10 
a = 8'd84; b = 8'd50;  #10 
a = 8'd84; b = 8'd51;  #10 
a = 8'd84; b = 8'd52;  #10 
a = 8'd84; b = 8'd53;  #10 
a = 8'd84; b = 8'd54;  #10 
a = 8'd84; b = 8'd55;  #10 
a = 8'd84; b = 8'd56;  #10 
a = 8'd84; b = 8'd57;  #10 
a = 8'd84; b = 8'd58;  #10 
a = 8'd84; b = 8'd59;  #10 
a = 8'd84; b = 8'd60;  #10 
a = 8'd84; b = 8'd61;  #10 
a = 8'd84; b = 8'd62;  #10 
a = 8'd84; b = 8'd63;  #10 
a = 8'd84; b = 8'd64;  #10 
a = 8'd84; b = 8'd65;  #10 
a = 8'd84; b = 8'd66;  #10 
a = 8'd84; b = 8'd67;  #10 
a = 8'd84; b = 8'd68;  #10 
a = 8'd84; b = 8'd69;  #10 
a = 8'd84; b = 8'd70;  #10 
a = 8'd84; b = 8'd71;  #10 
a = 8'd84; b = 8'd72;  #10 
a = 8'd84; b = 8'd73;  #10 
a = 8'd84; b = 8'd74;  #10 
a = 8'd84; b = 8'd75;  #10 
a = 8'd84; b = 8'd76;  #10 
a = 8'd84; b = 8'd77;  #10 
a = 8'd84; b = 8'd78;  #10 
a = 8'd84; b = 8'd79;  #10 
a = 8'd84; b = 8'd80;  #10 
a = 8'd84; b = 8'd81;  #10 
a = 8'd84; b = 8'd82;  #10 
a = 8'd84; b = 8'd83;  #10 
a = 8'd84; b = 8'd84;  #10 
a = 8'd84; b = 8'd85;  #10 
a = 8'd84; b = 8'd86;  #10 
a = 8'd84; b = 8'd87;  #10 
a = 8'd84; b = 8'd88;  #10 
a = 8'd84; b = 8'd89;  #10 
a = 8'd84; b = 8'd90;  #10 
a = 8'd84; b = 8'd91;  #10 
a = 8'd84; b = 8'd92;  #10 
a = 8'd84; b = 8'd93;  #10 
a = 8'd84; b = 8'd94;  #10 
a = 8'd84; b = 8'd95;  #10 
a = 8'd84; b = 8'd96;  #10 
a = 8'd84; b = 8'd97;  #10 
a = 8'd84; b = 8'd98;  #10 
a = 8'd84; b = 8'd99;  #10 
a = 8'd84; b = 8'd100;  #10 
a = 8'd84; b = 8'd101;  #10 
a = 8'd84; b = 8'd102;  #10 
a = 8'd84; b = 8'd103;  #10 
a = 8'd84; b = 8'd104;  #10 
a = 8'd84; b = 8'd105;  #10 
a = 8'd84; b = 8'd106;  #10 
a = 8'd84; b = 8'd107;  #10 
a = 8'd84; b = 8'd108;  #10 
a = 8'd84; b = 8'd109;  #10 
a = 8'd84; b = 8'd110;  #10 
a = 8'd84; b = 8'd111;  #10 
a = 8'd84; b = 8'd112;  #10 
a = 8'd84; b = 8'd113;  #10 
a = 8'd84; b = 8'd114;  #10 
a = 8'd84; b = 8'd115;  #10 
a = 8'd84; b = 8'd116;  #10 
a = 8'd84; b = 8'd117;  #10 
a = 8'd84; b = 8'd118;  #10 
a = 8'd84; b = 8'd119;  #10 
a = 8'd84; b = 8'd120;  #10 
a = 8'd84; b = 8'd121;  #10 
a = 8'd84; b = 8'd122;  #10 
a = 8'd84; b = 8'd123;  #10 
a = 8'd84; b = 8'd124;  #10 
a = 8'd84; b = 8'd125;  #10 
a = 8'd84; b = 8'd126;  #10 
a = 8'd84; b = 8'd127;  #10 
a = 8'd84; b = 8'd128;  #10 
a = 8'd84; b = 8'd129;  #10 
a = 8'd84; b = 8'd130;  #10 
a = 8'd84; b = 8'd131;  #10 
a = 8'd84; b = 8'd132;  #10 
a = 8'd84; b = 8'd133;  #10 
a = 8'd84; b = 8'd134;  #10 
a = 8'd84; b = 8'd135;  #10 
a = 8'd84; b = 8'd136;  #10 
a = 8'd84; b = 8'd137;  #10 
a = 8'd84; b = 8'd138;  #10 
a = 8'd84; b = 8'd139;  #10 
a = 8'd84; b = 8'd140;  #10 
a = 8'd84; b = 8'd141;  #10 
a = 8'd84; b = 8'd142;  #10 
a = 8'd84; b = 8'd143;  #10 
a = 8'd84; b = 8'd144;  #10 
a = 8'd84; b = 8'd145;  #10 
a = 8'd84; b = 8'd146;  #10 
a = 8'd84; b = 8'd147;  #10 
a = 8'd84; b = 8'd148;  #10 
a = 8'd84; b = 8'd149;  #10 
a = 8'd84; b = 8'd150;  #10 
a = 8'd84; b = 8'd151;  #10 
a = 8'd84; b = 8'd152;  #10 
a = 8'd84; b = 8'd153;  #10 
a = 8'd84; b = 8'd154;  #10 
a = 8'd84; b = 8'd155;  #10 
a = 8'd84; b = 8'd156;  #10 
a = 8'd84; b = 8'd157;  #10 
a = 8'd84; b = 8'd158;  #10 
a = 8'd84; b = 8'd159;  #10 
a = 8'd84; b = 8'd160;  #10 
a = 8'd84; b = 8'd161;  #10 
a = 8'd84; b = 8'd162;  #10 
a = 8'd84; b = 8'd163;  #10 
a = 8'd84; b = 8'd164;  #10 
a = 8'd84; b = 8'd165;  #10 
a = 8'd84; b = 8'd166;  #10 
a = 8'd84; b = 8'd167;  #10 
a = 8'd84; b = 8'd168;  #10 
a = 8'd84; b = 8'd169;  #10 
a = 8'd84; b = 8'd170;  #10 
a = 8'd84; b = 8'd171;  #10 
a = 8'd84; b = 8'd172;  #10 
a = 8'd84; b = 8'd173;  #10 
a = 8'd84; b = 8'd174;  #10 
a = 8'd84; b = 8'd175;  #10 
a = 8'd84; b = 8'd176;  #10 
a = 8'd84; b = 8'd177;  #10 
a = 8'd84; b = 8'd178;  #10 
a = 8'd84; b = 8'd179;  #10 
a = 8'd84; b = 8'd180;  #10 
a = 8'd84; b = 8'd181;  #10 
a = 8'd84; b = 8'd182;  #10 
a = 8'd84; b = 8'd183;  #10 
a = 8'd84; b = 8'd184;  #10 
a = 8'd84; b = 8'd185;  #10 
a = 8'd84; b = 8'd186;  #10 
a = 8'd84; b = 8'd187;  #10 
a = 8'd84; b = 8'd188;  #10 
a = 8'd84; b = 8'd189;  #10 
a = 8'd84; b = 8'd190;  #10 
a = 8'd84; b = 8'd191;  #10 
a = 8'd84; b = 8'd192;  #10 
a = 8'd84; b = 8'd193;  #10 
a = 8'd84; b = 8'd194;  #10 
a = 8'd84; b = 8'd195;  #10 
a = 8'd84; b = 8'd196;  #10 
a = 8'd84; b = 8'd197;  #10 
a = 8'd84; b = 8'd198;  #10 
a = 8'd84; b = 8'd199;  #10 
a = 8'd84; b = 8'd200;  #10 
a = 8'd84; b = 8'd201;  #10 
a = 8'd84; b = 8'd202;  #10 
a = 8'd84; b = 8'd203;  #10 
a = 8'd84; b = 8'd204;  #10 
a = 8'd84; b = 8'd205;  #10 
a = 8'd84; b = 8'd206;  #10 
a = 8'd84; b = 8'd207;  #10 
a = 8'd84; b = 8'd208;  #10 
a = 8'd84; b = 8'd209;  #10 
a = 8'd84; b = 8'd210;  #10 
a = 8'd84; b = 8'd211;  #10 
a = 8'd84; b = 8'd212;  #10 
a = 8'd84; b = 8'd213;  #10 
a = 8'd84; b = 8'd214;  #10 
a = 8'd84; b = 8'd215;  #10 
a = 8'd84; b = 8'd216;  #10 
a = 8'd84; b = 8'd217;  #10 
a = 8'd84; b = 8'd218;  #10 
a = 8'd84; b = 8'd219;  #10 
a = 8'd84; b = 8'd220;  #10 
a = 8'd84; b = 8'd221;  #10 
a = 8'd84; b = 8'd222;  #10 
a = 8'd84; b = 8'd223;  #10 
a = 8'd84; b = 8'd224;  #10 
a = 8'd84; b = 8'd225;  #10 
a = 8'd84; b = 8'd226;  #10 
a = 8'd84; b = 8'd227;  #10 
a = 8'd84; b = 8'd228;  #10 
a = 8'd84; b = 8'd229;  #10 
a = 8'd84; b = 8'd230;  #10 
a = 8'd84; b = 8'd231;  #10 
a = 8'd84; b = 8'd232;  #10 
a = 8'd84; b = 8'd233;  #10 
a = 8'd84; b = 8'd234;  #10 
a = 8'd84; b = 8'd235;  #10 
a = 8'd84; b = 8'd236;  #10 
a = 8'd84; b = 8'd237;  #10 
a = 8'd84; b = 8'd238;  #10 
a = 8'd84; b = 8'd239;  #10 
a = 8'd84; b = 8'd240;  #10 
a = 8'd84; b = 8'd241;  #10 
a = 8'd84; b = 8'd242;  #10 
a = 8'd84; b = 8'd243;  #10 
a = 8'd84; b = 8'd244;  #10 
a = 8'd84; b = 8'd245;  #10 
a = 8'd84; b = 8'd246;  #10 
a = 8'd84; b = 8'd247;  #10 
a = 8'd84; b = 8'd248;  #10 
a = 8'd84; b = 8'd249;  #10 
a = 8'd84; b = 8'd250;  #10 
a = 8'd84; b = 8'd251;  #10 
a = 8'd84; b = 8'd252;  #10 
a = 8'd84; b = 8'd253;  #10 
a = 8'd84; b = 8'd254;  #10 
a = 8'd84; b = 8'd255;  #10 
a = 8'd85; b = 8'd0;  #10 
a = 8'd85; b = 8'd1;  #10 
a = 8'd85; b = 8'd2;  #10 
a = 8'd85; b = 8'd3;  #10 
a = 8'd85; b = 8'd4;  #10 
a = 8'd85; b = 8'd5;  #10 
a = 8'd85; b = 8'd6;  #10 
a = 8'd85; b = 8'd7;  #10 
a = 8'd85; b = 8'd8;  #10 
a = 8'd85; b = 8'd9;  #10 
a = 8'd85; b = 8'd10;  #10 
a = 8'd85; b = 8'd11;  #10 
a = 8'd85; b = 8'd12;  #10 
a = 8'd85; b = 8'd13;  #10 
a = 8'd85; b = 8'd14;  #10 
a = 8'd85; b = 8'd15;  #10 
a = 8'd85; b = 8'd16;  #10 
a = 8'd85; b = 8'd17;  #10 
a = 8'd85; b = 8'd18;  #10 
a = 8'd85; b = 8'd19;  #10 
a = 8'd85; b = 8'd20;  #10 
a = 8'd85; b = 8'd21;  #10 
a = 8'd85; b = 8'd22;  #10 
a = 8'd85; b = 8'd23;  #10 
a = 8'd85; b = 8'd24;  #10 
a = 8'd85; b = 8'd25;  #10 
a = 8'd85; b = 8'd26;  #10 
a = 8'd85; b = 8'd27;  #10 
a = 8'd85; b = 8'd28;  #10 
a = 8'd85; b = 8'd29;  #10 
a = 8'd85; b = 8'd30;  #10 
a = 8'd85; b = 8'd31;  #10 
a = 8'd85; b = 8'd32;  #10 
a = 8'd85; b = 8'd33;  #10 
a = 8'd85; b = 8'd34;  #10 
a = 8'd85; b = 8'd35;  #10 
a = 8'd85; b = 8'd36;  #10 
a = 8'd85; b = 8'd37;  #10 
a = 8'd85; b = 8'd38;  #10 
a = 8'd85; b = 8'd39;  #10 
a = 8'd85; b = 8'd40;  #10 
a = 8'd85; b = 8'd41;  #10 
a = 8'd85; b = 8'd42;  #10 
a = 8'd85; b = 8'd43;  #10 
a = 8'd85; b = 8'd44;  #10 
a = 8'd85; b = 8'd45;  #10 
a = 8'd85; b = 8'd46;  #10 
a = 8'd85; b = 8'd47;  #10 
a = 8'd85; b = 8'd48;  #10 
a = 8'd85; b = 8'd49;  #10 
a = 8'd85; b = 8'd50;  #10 
a = 8'd85; b = 8'd51;  #10 
a = 8'd85; b = 8'd52;  #10 
a = 8'd85; b = 8'd53;  #10 
a = 8'd85; b = 8'd54;  #10 
a = 8'd85; b = 8'd55;  #10 
a = 8'd85; b = 8'd56;  #10 
a = 8'd85; b = 8'd57;  #10 
a = 8'd85; b = 8'd58;  #10 
a = 8'd85; b = 8'd59;  #10 
a = 8'd85; b = 8'd60;  #10 
a = 8'd85; b = 8'd61;  #10 
a = 8'd85; b = 8'd62;  #10 
a = 8'd85; b = 8'd63;  #10 
a = 8'd85; b = 8'd64;  #10 
a = 8'd85; b = 8'd65;  #10 
a = 8'd85; b = 8'd66;  #10 
a = 8'd85; b = 8'd67;  #10 
a = 8'd85; b = 8'd68;  #10 
a = 8'd85; b = 8'd69;  #10 
a = 8'd85; b = 8'd70;  #10 
a = 8'd85; b = 8'd71;  #10 
a = 8'd85; b = 8'd72;  #10 
a = 8'd85; b = 8'd73;  #10 
a = 8'd85; b = 8'd74;  #10 
a = 8'd85; b = 8'd75;  #10 
a = 8'd85; b = 8'd76;  #10 
a = 8'd85; b = 8'd77;  #10 
a = 8'd85; b = 8'd78;  #10 
a = 8'd85; b = 8'd79;  #10 
a = 8'd85; b = 8'd80;  #10 
a = 8'd85; b = 8'd81;  #10 
a = 8'd85; b = 8'd82;  #10 
a = 8'd85; b = 8'd83;  #10 
a = 8'd85; b = 8'd84;  #10 
a = 8'd85; b = 8'd85;  #10 
a = 8'd85; b = 8'd86;  #10 
a = 8'd85; b = 8'd87;  #10 
a = 8'd85; b = 8'd88;  #10 
a = 8'd85; b = 8'd89;  #10 
a = 8'd85; b = 8'd90;  #10 
a = 8'd85; b = 8'd91;  #10 
a = 8'd85; b = 8'd92;  #10 
a = 8'd85; b = 8'd93;  #10 
a = 8'd85; b = 8'd94;  #10 
a = 8'd85; b = 8'd95;  #10 
a = 8'd85; b = 8'd96;  #10 
a = 8'd85; b = 8'd97;  #10 
a = 8'd85; b = 8'd98;  #10 
a = 8'd85; b = 8'd99;  #10 
a = 8'd85; b = 8'd100;  #10 
a = 8'd85; b = 8'd101;  #10 
a = 8'd85; b = 8'd102;  #10 
a = 8'd85; b = 8'd103;  #10 
a = 8'd85; b = 8'd104;  #10 
a = 8'd85; b = 8'd105;  #10 
a = 8'd85; b = 8'd106;  #10 
a = 8'd85; b = 8'd107;  #10 
a = 8'd85; b = 8'd108;  #10 
a = 8'd85; b = 8'd109;  #10 
a = 8'd85; b = 8'd110;  #10 
a = 8'd85; b = 8'd111;  #10 
a = 8'd85; b = 8'd112;  #10 
a = 8'd85; b = 8'd113;  #10 
a = 8'd85; b = 8'd114;  #10 
a = 8'd85; b = 8'd115;  #10 
a = 8'd85; b = 8'd116;  #10 
a = 8'd85; b = 8'd117;  #10 
a = 8'd85; b = 8'd118;  #10 
a = 8'd85; b = 8'd119;  #10 
a = 8'd85; b = 8'd120;  #10 
a = 8'd85; b = 8'd121;  #10 
a = 8'd85; b = 8'd122;  #10 
a = 8'd85; b = 8'd123;  #10 
a = 8'd85; b = 8'd124;  #10 
a = 8'd85; b = 8'd125;  #10 
a = 8'd85; b = 8'd126;  #10 
a = 8'd85; b = 8'd127;  #10 
a = 8'd85; b = 8'd128;  #10 
a = 8'd85; b = 8'd129;  #10 
a = 8'd85; b = 8'd130;  #10 
a = 8'd85; b = 8'd131;  #10 
a = 8'd85; b = 8'd132;  #10 
a = 8'd85; b = 8'd133;  #10 
a = 8'd85; b = 8'd134;  #10 
a = 8'd85; b = 8'd135;  #10 
a = 8'd85; b = 8'd136;  #10 
a = 8'd85; b = 8'd137;  #10 
a = 8'd85; b = 8'd138;  #10 
a = 8'd85; b = 8'd139;  #10 
a = 8'd85; b = 8'd140;  #10 
a = 8'd85; b = 8'd141;  #10 
a = 8'd85; b = 8'd142;  #10 
a = 8'd85; b = 8'd143;  #10 
a = 8'd85; b = 8'd144;  #10 
a = 8'd85; b = 8'd145;  #10 
a = 8'd85; b = 8'd146;  #10 
a = 8'd85; b = 8'd147;  #10 
a = 8'd85; b = 8'd148;  #10 
a = 8'd85; b = 8'd149;  #10 
a = 8'd85; b = 8'd150;  #10 
a = 8'd85; b = 8'd151;  #10 
a = 8'd85; b = 8'd152;  #10 
a = 8'd85; b = 8'd153;  #10 
a = 8'd85; b = 8'd154;  #10 
a = 8'd85; b = 8'd155;  #10 
a = 8'd85; b = 8'd156;  #10 
a = 8'd85; b = 8'd157;  #10 
a = 8'd85; b = 8'd158;  #10 
a = 8'd85; b = 8'd159;  #10 
a = 8'd85; b = 8'd160;  #10 
a = 8'd85; b = 8'd161;  #10 
a = 8'd85; b = 8'd162;  #10 
a = 8'd85; b = 8'd163;  #10 
a = 8'd85; b = 8'd164;  #10 
a = 8'd85; b = 8'd165;  #10 
a = 8'd85; b = 8'd166;  #10 
a = 8'd85; b = 8'd167;  #10 
a = 8'd85; b = 8'd168;  #10 
a = 8'd85; b = 8'd169;  #10 
a = 8'd85; b = 8'd170;  #10 
a = 8'd85; b = 8'd171;  #10 
a = 8'd85; b = 8'd172;  #10 
a = 8'd85; b = 8'd173;  #10 
a = 8'd85; b = 8'd174;  #10 
a = 8'd85; b = 8'd175;  #10 
a = 8'd85; b = 8'd176;  #10 
a = 8'd85; b = 8'd177;  #10 
a = 8'd85; b = 8'd178;  #10 
a = 8'd85; b = 8'd179;  #10 
a = 8'd85; b = 8'd180;  #10 
a = 8'd85; b = 8'd181;  #10 
a = 8'd85; b = 8'd182;  #10 
a = 8'd85; b = 8'd183;  #10 
a = 8'd85; b = 8'd184;  #10 
a = 8'd85; b = 8'd185;  #10 
a = 8'd85; b = 8'd186;  #10 
a = 8'd85; b = 8'd187;  #10 
a = 8'd85; b = 8'd188;  #10 
a = 8'd85; b = 8'd189;  #10 
a = 8'd85; b = 8'd190;  #10 
a = 8'd85; b = 8'd191;  #10 
a = 8'd85; b = 8'd192;  #10 
a = 8'd85; b = 8'd193;  #10 
a = 8'd85; b = 8'd194;  #10 
a = 8'd85; b = 8'd195;  #10 
a = 8'd85; b = 8'd196;  #10 
a = 8'd85; b = 8'd197;  #10 
a = 8'd85; b = 8'd198;  #10 
a = 8'd85; b = 8'd199;  #10 
a = 8'd85; b = 8'd200;  #10 
a = 8'd85; b = 8'd201;  #10 
a = 8'd85; b = 8'd202;  #10 
a = 8'd85; b = 8'd203;  #10 
a = 8'd85; b = 8'd204;  #10 
a = 8'd85; b = 8'd205;  #10 
a = 8'd85; b = 8'd206;  #10 
a = 8'd85; b = 8'd207;  #10 
a = 8'd85; b = 8'd208;  #10 
a = 8'd85; b = 8'd209;  #10 
a = 8'd85; b = 8'd210;  #10 
a = 8'd85; b = 8'd211;  #10 
a = 8'd85; b = 8'd212;  #10 
a = 8'd85; b = 8'd213;  #10 
a = 8'd85; b = 8'd214;  #10 
a = 8'd85; b = 8'd215;  #10 
a = 8'd85; b = 8'd216;  #10 
a = 8'd85; b = 8'd217;  #10 
a = 8'd85; b = 8'd218;  #10 
a = 8'd85; b = 8'd219;  #10 
a = 8'd85; b = 8'd220;  #10 
a = 8'd85; b = 8'd221;  #10 
a = 8'd85; b = 8'd222;  #10 
a = 8'd85; b = 8'd223;  #10 
a = 8'd85; b = 8'd224;  #10 
a = 8'd85; b = 8'd225;  #10 
a = 8'd85; b = 8'd226;  #10 
a = 8'd85; b = 8'd227;  #10 
a = 8'd85; b = 8'd228;  #10 
a = 8'd85; b = 8'd229;  #10 
a = 8'd85; b = 8'd230;  #10 
a = 8'd85; b = 8'd231;  #10 
a = 8'd85; b = 8'd232;  #10 
a = 8'd85; b = 8'd233;  #10 
a = 8'd85; b = 8'd234;  #10 
a = 8'd85; b = 8'd235;  #10 
a = 8'd85; b = 8'd236;  #10 
a = 8'd85; b = 8'd237;  #10 
a = 8'd85; b = 8'd238;  #10 
a = 8'd85; b = 8'd239;  #10 
a = 8'd85; b = 8'd240;  #10 
a = 8'd85; b = 8'd241;  #10 
a = 8'd85; b = 8'd242;  #10 
a = 8'd85; b = 8'd243;  #10 
a = 8'd85; b = 8'd244;  #10 
a = 8'd85; b = 8'd245;  #10 
a = 8'd85; b = 8'd246;  #10 
a = 8'd85; b = 8'd247;  #10 
a = 8'd85; b = 8'd248;  #10 
a = 8'd85; b = 8'd249;  #10 
a = 8'd85; b = 8'd250;  #10 
a = 8'd85; b = 8'd251;  #10 
a = 8'd85; b = 8'd252;  #10 
a = 8'd85; b = 8'd253;  #10 
a = 8'd85; b = 8'd254;  #10 
a = 8'd85; b = 8'd255;  #10 
a = 8'd86; b = 8'd0;  #10 
a = 8'd86; b = 8'd1;  #10 
a = 8'd86; b = 8'd2;  #10 
a = 8'd86; b = 8'd3;  #10 
a = 8'd86; b = 8'd4;  #10 
a = 8'd86; b = 8'd5;  #10 
a = 8'd86; b = 8'd6;  #10 
a = 8'd86; b = 8'd7;  #10 
a = 8'd86; b = 8'd8;  #10 
a = 8'd86; b = 8'd9;  #10 
a = 8'd86; b = 8'd10;  #10 
a = 8'd86; b = 8'd11;  #10 
a = 8'd86; b = 8'd12;  #10 
a = 8'd86; b = 8'd13;  #10 
a = 8'd86; b = 8'd14;  #10 
a = 8'd86; b = 8'd15;  #10 
a = 8'd86; b = 8'd16;  #10 
a = 8'd86; b = 8'd17;  #10 
a = 8'd86; b = 8'd18;  #10 
a = 8'd86; b = 8'd19;  #10 
a = 8'd86; b = 8'd20;  #10 
a = 8'd86; b = 8'd21;  #10 
a = 8'd86; b = 8'd22;  #10 
a = 8'd86; b = 8'd23;  #10 
a = 8'd86; b = 8'd24;  #10 
a = 8'd86; b = 8'd25;  #10 
a = 8'd86; b = 8'd26;  #10 
a = 8'd86; b = 8'd27;  #10 
a = 8'd86; b = 8'd28;  #10 
a = 8'd86; b = 8'd29;  #10 
a = 8'd86; b = 8'd30;  #10 
a = 8'd86; b = 8'd31;  #10 
a = 8'd86; b = 8'd32;  #10 
a = 8'd86; b = 8'd33;  #10 
a = 8'd86; b = 8'd34;  #10 
a = 8'd86; b = 8'd35;  #10 
a = 8'd86; b = 8'd36;  #10 
a = 8'd86; b = 8'd37;  #10 
a = 8'd86; b = 8'd38;  #10 
a = 8'd86; b = 8'd39;  #10 
a = 8'd86; b = 8'd40;  #10 
a = 8'd86; b = 8'd41;  #10 
a = 8'd86; b = 8'd42;  #10 
a = 8'd86; b = 8'd43;  #10 
a = 8'd86; b = 8'd44;  #10 
a = 8'd86; b = 8'd45;  #10 
a = 8'd86; b = 8'd46;  #10 
a = 8'd86; b = 8'd47;  #10 
a = 8'd86; b = 8'd48;  #10 
a = 8'd86; b = 8'd49;  #10 
a = 8'd86; b = 8'd50;  #10 
a = 8'd86; b = 8'd51;  #10 
a = 8'd86; b = 8'd52;  #10 
a = 8'd86; b = 8'd53;  #10 
a = 8'd86; b = 8'd54;  #10 
a = 8'd86; b = 8'd55;  #10 
a = 8'd86; b = 8'd56;  #10 
a = 8'd86; b = 8'd57;  #10 
a = 8'd86; b = 8'd58;  #10 
a = 8'd86; b = 8'd59;  #10 
a = 8'd86; b = 8'd60;  #10 
a = 8'd86; b = 8'd61;  #10 
a = 8'd86; b = 8'd62;  #10 
a = 8'd86; b = 8'd63;  #10 
a = 8'd86; b = 8'd64;  #10 
a = 8'd86; b = 8'd65;  #10 
a = 8'd86; b = 8'd66;  #10 
a = 8'd86; b = 8'd67;  #10 
a = 8'd86; b = 8'd68;  #10 
a = 8'd86; b = 8'd69;  #10 
a = 8'd86; b = 8'd70;  #10 
a = 8'd86; b = 8'd71;  #10 
a = 8'd86; b = 8'd72;  #10 
a = 8'd86; b = 8'd73;  #10 
a = 8'd86; b = 8'd74;  #10 
a = 8'd86; b = 8'd75;  #10 
a = 8'd86; b = 8'd76;  #10 
a = 8'd86; b = 8'd77;  #10 
a = 8'd86; b = 8'd78;  #10 
a = 8'd86; b = 8'd79;  #10 
a = 8'd86; b = 8'd80;  #10 
a = 8'd86; b = 8'd81;  #10 
a = 8'd86; b = 8'd82;  #10 
a = 8'd86; b = 8'd83;  #10 
a = 8'd86; b = 8'd84;  #10 
a = 8'd86; b = 8'd85;  #10 
a = 8'd86; b = 8'd86;  #10 
a = 8'd86; b = 8'd87;  #10 
a = 8'd86; b = 8'd88;  #10 
a = 8'd86; b = 8'd89;  #10 
a = 8'd86; b = 8'd90;  #10 
a = 8'd86; b = 8'd91;  #10 
a = 8'd86; b = 8'd92;  #10 
a = 8'd86; b = 8'd93;  #10 
a = 8'd86; b = 8'd94;  #10 
a = 8'd86; b = 8'd95;  #10 
a = 8'd86; b = 8'd96;  #10 
a = 8'd86; b = 8'd97;  #10 
a = 8'd86; b = 8'd98;  #10 
a = 8'd86; b = 8'd99;  #10 
a = 8'd86; b = 8'd100;  #10 
a = 8'd86; b = 8'd101;  #10 
a = 8'd86; b = 8'd102;  #10 
a = 8'd86; b = 8'd103;  #10 
a = 8'd86; b = 8'd104;  #10 
a = 8'd86; b = 8'd105;  #10 
a = 8'd86; b = 8'd106;  #10 
a = 8'd86; b = 8'd107;  #10 
a = 8'd86; b = 8'd108;  #10 
a = 8'd86; b = 8'd109;  #10 
a = 8'd86; b = 8'd110;  #10 
a = 8'd86; b = 8'd111;  #10 
a = 8'd86; b = 8'd112;  #10 
a = 8'd86; b = 8'd113;  #10 
a = 8'd86; b = 8'd114;  #10 
a = 8'd86; b = 8'd115;  #10 
a = 8'd86; b = 8'd116;  #10 
a = 8'd86; b = 8'd117;  #10 
a = 8'd86; b = 8'd118;  #10 
a = 8'd86; b = 8'd119;  #10 
a = 8'd86; b = 8'd120;  #10 
a = 8'd86; b = 8'd121;  #10 
a = 8'd86; b = 8'd122;  #10 
a = 8'd86; b = 8'd123;  #10 
a = 8'd86; b = 8'd124;  #10 
a = 8'd86; b = 8'd125;  #10 
a = 8'd86; b = 8'd126;  #10 
a = 8'd86; b = 8'd127;  #10 
a = 8'd86; b = 8'd128;  #10 
a = 8'd86; b = 8'd129;  #10 
a = 8'd86; b = 8'd130;  #10 
a = 8'd86; b = 8'd131;  #10 
a = 8'd86; b = 8'd132;  #10 
a = 8'd86; b = 8'd133;  #10 
a = 8'd86; b = 8'd134;  #10 
a = 8'd86; b = 8'd135;  #10 
a = 8'd86; b = 8'd136;  #10 
a = 8'd86; b = 8'd137;  #10 
a = 8'd86; b = 8'd138;  #10 
a = 8'd86; b = 8'd139;  #10 
a = 8'd86; b = 8'd140;  #10 
a = 8'd86; b = 8'd141;  #10 
a = 8'd86; b = 8'd142;  #10 
a = 8'd86; b = 8'd143;  #10 
a = 8'd86; b = 8'd144;  #10 
a = 8'd86; b = 8'd145;  #10 
a = 8'd86; b = 8'd146;  #10 
a = 8'd86; b = 8'd147;  #10 
a = 8'd86; b = 8'd148;  #10 
a = 8'd86; b = 8'd149;  #10 
a = 8'd86; b = 8'd150;  #10 
a = 8'd86; b = 8'd151;  #10 
a = 8'd86; b = 8'd152;  #10 
a = 8'd86; b = 8'd153;  #10 
a = 8'd86; b = 8'd154;  #10 
a = 8'd86; b = 8'd155;  #10 
a = 8'd86; b = 8'd156;  #10 
a = 8'd86; b = 8'd157;  #10 
a = 8'd86; b = 8'd158;  #10 
a = 8'd86; b = 8'd159;  #10 
a = 8'd86; b = 8'd160;  #10 
a = 8'd86; b = 8'd161;  #10 
a = 8'd86; b = 8'd162;  #10 
a = 8'd86; b = 8'd163;  #10 
a = 8'd86; b = 8'd164;  #10 
a = 8'd86; b = 8'd165;  #10 
a = 8'd86; b = 8'd166;  #10 
a = 8'd86; b = 8'd167;  #10 
a = 8'd86; b = 8'd168;  #10 
a = 8'd86; b = 8'd169;  #10 
a = 8'd86; b = 8'd170;  #10 
a = 8'd86; b = 8'd171;  #10 
a = 8'd86; b = 8'd172;  #10 
a = 8'd86; b = 8'd173;  #10 
a = 8'd86; b = 8'd174;  #10 
a = 8'd86; b = 8'd175;  #10 
a = 8'd86; b = 8'd176;  #10 
a = 8'd86; b = 8'd177;  #10 
a = 8'd86; b = 8'd178;  #10 
a = 8'd86; b = 8'd179;  #10 
a = 8'd86; b = 8'd180;  #10 
a = 8'd86; b = 8'd181;  #10 
a = 8'd86; b = 8'd182;  #10 
a = 8'd86; b = 8'd183;  #10 
a = 8'd86; b = 8'd184;  #10 
a = 8'd86; b = 8'd185;  #10 
a = 8'd86; b = 8'd186;  #10 
a = 8'd86; b = 8'd187;  #10 
a = 8'd86; b = 8'd188;  #10 
a = 8'd86; b = 8'd189;  #10 
a = 8'd86; b = 8'd190;  #10 
a = 8'd86; b = 8'd191;  #10 
a = 8'd86; b = 8'd192;  #10 
a = 8'd86; b = 8'd193;  #10 
a = 8'd86; b = 8'd194;  #10 
a = 8'd86; b = 8'd195;  #10 
a = 8'd86; b = 8'd196;  #10 
a = 8'd86; b = 8'd197;  #10 
a = 8'd86; b = 8'd198;  #10 
a = 8'd86; b = 8'd199;  #10 
a = 8'd86; b = 8'd200;  #10 
a = 8'd86; b = 8'd201;  #10 
a = 8'd86; b = 8'd202;  #10 
a = 8'd86; b = 8'd203;  #10 
a = 8'd86; b = 8'd204;  #10 
a = 8'd86; b = 8'd205;  #10 
a = 8'd86; b = 8'd206;  #10 
a = 8'd86; b = 8'd207;  #10 
a = 8'd86; b = 8'd208;  #10 
a = 8'd86; b = 8'd209;  #10 
a = 8'd86; b = 8'd210;  #10 
a = 8'd86; b = 8'd211;  #10 
a = 8'd86; b = 8'd212;  #10 
a = 8'd86; b = 8'd213;  #10 
a = 8'd86; b = 8'd214;  #10 
a = 8'd86; b = 8'd215;  #10 
a = 8'd86; b = 8'd216;  #10 
a = 8'd86; b = 8'd217;  #10 
a = 8'd86; b = 8'd218;  #10 
a = 8'd86; b = 8'd219;  #10 
a = 8'd86; b = 8'd220;  #10 
a = 8'd86; b = 8'd221;  #10 
a = 8'd86; b = 8'd222;  #10 
a = 8'd86; b = 8'd223;  #10 
a = 8'd86; b = 8'd224;  #10 
a = 8'd86; b = 8'd225;  #10 
a = 8'd86; b = 8'd226;  #10 
a = 8'd86; b = 8'd227;  #10 
a = 8'd86; b = 8'd228;  #10 
a = 8'd86; b = 8'd229;  #10 
a = 8'd86; b = 8'd230;  #10 
a = 8'd86; b = 8'd231;  #10 
a = 8'd86; b = 8'd232;  #10 
a = 8'd86; b = 8'd233;  #10 
a = 8'd86; b = 8'd234;  #10 
a = 8'd86; b = 8'd235;  #10 
a = 8'd86; b = 8'd236;  #10 
a = 8'd86; b = 8'd237;  #10 
a = 8'd86; b = 8'd238;  #10 
a = 8'd86; b = 8'd239;  #10 
a = 8'd86; b = 8'd240;  #10 
a = 8'd86; b = 8'd241;  #10 
a = 8'd86; b = 8'd242;  #10 
a = 8'd86; b = 8'd243;  #10 
a = 8'd86; b = 8'd244;  #10 
a = 8'd86; b = 8'd245;  #10 
a = 8'd86; b = 8'd246;  #10 
a = 8'd86; b = 8'd247;  #10 
a = 8'd86; b = 8'd248;  #10 
a = 8'd86; b = 8'd249;  #10 
a = 8'd86; b = 8'd250;  #10 
a = 8'd86; b = 8'd251;  #10 
a = 8'd86; b = 8'd252;  #10 
a = 8'd86; b = 8'd253;  #10 
a = 8'd86; b = 8'd254;  #10 
a = 8'd86; b = 8'd255;  #10 
a = 8'd87; b = 8'd0;  #10 
a = 8'd87; b = 8'd1;  #10 
a = 8'd87; b = 8'd2;  #10 
a = 8'd87; b = 8'd3;  #10 
a = 8'd87; b = 8'd4;  #10 
a = 8'd87; b = 8'd5;  #10 
a = 8'd87; b = 8'd6;  #10 
a = 8'd87; b = 8'd7;  #10 
a = 8'd87; b = 8'd8;  #10 
a = 8'd87; b = 8'd9;  #10 
a = 8'd87; b = 8'd10;  #10 
a = 8'd87; b = 8'd11;  #10 
a = 8'd87; b = 8'd12;  #10 
a = 8'd87; b = 8'd13;  #10 
a = 8'd87; b = 8'd14;  #10 
a = 8'd87; b = 8'd15;  #10 
a = 8'd87; b = 8'd16;  #10 
a = 8'd87; b = 8'd17;  #10 
a = 8'd87; b = 8'd18;  #10 
a = 8'd87; b = 8'd19;  #10 
a = 8'd87; b = 8'd20;  #10 
a = 8'd87; b = 8'd21;  #10 
a = 8'd87; b = 8'd22;  #10 
a = 8'd87; b = 8'd23;  #10 
a = 8'd87; b = 8'd24;  #10 
a = 8'd87; b = 8'd25;  #10 
a = 8'd87; b = 8'd26;  #10 
a = 8'd87; b = 8'd27;  #10 
a = 8'd87; b = 8'd28;  #10 
a = 8'd87; b = 8'd29;  #10 
a = 8'd87; b = 8'd30;  #10 
a = 8'd87; b = 8'd31;  #10 
a = 8'd87; b = 8'd32;  #10 
a = 8'd87; b = 8'd33;  #10 
a = 8'd87; b = 8'd34;  #10 
a = 8'd87; b = 8'd35;  #10 
a = 8'd87; b = 8'd36;  #10 
a = 8'd87; b = 8'd37;  #10 
a = 8'd87; b = 8'd38;  #10 
a = 8'd87; b = 8'd39;  #10 
a = 8'd87; b = 8'd40;  #10 
a = 8'd87; b = 8'd41;  #10 
a = 8'd87; b = 8'd42;  #10 
a = 8'd87; b = 8'd43;  #10 
a = 8'd87; b = 8'd44;  #10 
a = 8'd87; b = 8'd45;  #10 
a = 8'd87; b = 8'd46;  #10 
a = 8'd87; b = 8'd47;  #10 
a = 8'd87; b = 8'd48;  #10 
a = 8'd87; b = 8'd49;  #10 
a = 8'd87; b = 8'd50;  #10 
a = 8'd87; b = 8'd51;  #10 
a = 8'd87; b = 8'd52;  #10 
a = 8'd87; b = 8'd53;  #10 
a = 8'd87; b = 8'd54;  #10 
a = 8'd87; b = 8'd55;  #10 
a = 8'd87; b = 8'd56;  #10 
a = 8'd87; b = 8'd57;  #10 
a = 8'd87; b = 8'd58;  #10 
a = 8'd87; b = 8'd59;  #10 
a = 8'd87; b = 8'd60;  #10 
a = 8'd87; b = 8'd61;  #10 
a = 8'd87; b = 8'd62;  #10 
a = 8'd87; b = 8'd63;  #10 
a = 8'd87; b = 8'd64;  #10 
a = 8'd87; b = 8'd65;  #10 
a = 8'd87; b = 8'd66;  #10 
a = 8'd87; b = 8'd67;  #10 
a = 8'd87; b = 8'd68;  #10 
a = 8'd87; b = 8'd69;  #10 
a = 8'd87; b = 8'd70;  #10 
a = 8'd87; b = 8'd71;  #10 
a = 8'd87; b = 8'd72;  #10 
a = 8'd87; b = 8'd73;  #10 
a = 8'd87; b = 8'd74;  #10 
a = 8'd87; b = 8'd75;  #10 
a = 8'd87; b = 8'd76;  #10 
a = 8'd87; b = 8'd77;  #10 
a = 8'd87; b = 8'd78;  #10 
a = 8'd87; b = 8'd79;  #10 
a = 8'd87; b = 8'd80;  #10 
a = 8'd87; b = 8'd81;  #10 
a = 8'd87; b = 8'd82;  #10 
a = 8'd87; b = 8'd83;  #10 
a = 8'd87; b = 8'd84;  #10 
a = 8'd87; b = 8'd85;  #10 
a = 8'd87; b = 8'd86;  #10 
a = 8'd87; b = 8'd87;  #10 
a = 8'd87; b = 8'd88;  #10 
a = 8'd87; b = 8'd89;  #10 
a = 8'd87; b = 8'd90;  #10 
a = 8'd87; b = 8'd91;  #10 
a = 8'd87; b = 8'd92;  #10 
a = 8'd87; b = 8'd93;  #10 
a = 8'd87; b = 8'd94;  #10 
a = 8'd87; b = 8'd95;  #10 
a = 8'd87; b = 8'd96;  #10 
a = 8'd87; b = 8'd97;  #10 
a = 8'd87; b = 8'd98;  #10 
a = 8'd87; b = 8'd99;  #10 
a = 8'd87; b = 8'd100;  #10 
a = 8'd87; b = 8'd101;  #10 
a = 8'd87; b = 8'd102;  #10 
a = 8'd87; b = 8'd103;  #10 
a = 8'd87; b = 8'd104;  #10 
a = 8'd87; b = 8'd105;  #10 
a = 8'd87; b = 8'd106;  #10 
a = 8'd87; b = 8'd107;  #10 
a = 8'd87; b = 8'd108;  #10 
a = 8'd87; b = 8'd109;  #10 
a = 8'd87; b = 8'd110;  #10 
a = 8'd87; b = 8'd111;  #10 
a = 8'd87; b = 8'd112;  #10 
a = 8'd87; b = 8'd113;  #10 
a = 8'd87; b = 8'd114;  #10 
a = 8'd87; b = 8'd115;  #10 
a = 8'd87; b = 8'd116;  #10 
a = 8'd87; b = 8'd117;  #10 
a = 8'd87; b = 8'd118;  #10 
a = 8'd87; b = 8'd119;  #10 
a = 8'd87; b = 8'd120;  #10 
a = 8'd87; b = 8'd121;  #10 
a = 8'd87; b = 8'd122;  #10 
a = 8'd87; b = 8'd123;  #10 
a = 8'd87; b = 8'd124;  #10 
a = 8'd87; b = 8'd125;  #10 
a = 8'd87; b = 8'd126;  #10 
a = 8'd87; b = 8'd127;  #10 
a = 8'd87; b = 8'd128;  #10 
a = 8'd87; b = 8'd129;  #10 
a = 8'd87; b = 8'd130;  #10 
a = 8'd87; b = 8'd131;  #10 
a = 8'd87; b = 8'd132;  #10 
a = 8'd87; b = 8'd133;  #10 
a = 8'd87; b = 8'd134;  #10 
a = 8'd87; b = 8'd135;  #10 
a = 8'd87; b = 8'd136;  #10 
a = 8'd87; b = 8'd137;  #10 
a = 8'd87; b = 8'd138;  #10 
a = 8'd87; b = 8'd139;  #10 
a = 8'd87; b = 8'd140;  #10 
a = 8'd87; b = 8'd141;  #10 
a = 8'd87; b = 8'd142;  #10 
a = 8'd87; b = 8'd143;  #10 
a = 8'd87; b = 8'd144;  #10 
a = 8'd87; b = 8'd145;  #10 
a = 8'd87; b = 8'd146;  #10 
a = 8'd87; b = 8'd147;  #10 
a = 8'd87; b = 8'd148;  #10 
a = 8'd87; b = 8'd149;  #10 
a = 8'd87; b = 8'd150;  #10 
a = 8'd87; b = 8'd151;  #10 
a = 8'd87; b = 8'd152;  #10 
a = 8'd87; b = 8'd153;  #10 
a = 8'd87; b = 8'd154;  #10 
a = 8'd87; b = 8'd155;  #10 
a = 8'd87; b = 8'd156;  #10 
a = 8'd87; b = 8'd157;  #10 
a = 8'd87; b = 8'd158;  #10 
a = 8'd87; b = 8'd159;  #10 
a = 8'd87; b = 8'd160;  #10 
a = 8'd87; b = 8'd161;  #10 
a = 8'd87; b = 8'd162;  #10 
a = 8'd87; b = 8'd163;  #10 
a = 8'd87; b = 8'd164;  #10 
a = 8'd87; b = 8'd165;  #10 
a = 8'd87; b = 8'd166;  #10 
a = 8'd87; b = 8'd167;  #10 
a = 8'd87; b = 8'd168;  #10 
a = 8'd87; b = 8'd169;  #10 
a = 8'd87; b = 8'd170;  #10 
a = 8'd87; b = 8'd171;  #10 
a = 8'd87; b = 8'd172;  #10 
a = 8'd87; b = 8'd173;  #10 
a = 8'd87; b = 8'd174;  #10 
a = 8'd87; b = 8'd175;  #10 
a = 8'd87; b = 8'd176;  #10 
a = 8'd87; b = 8'd177;  #10 
a = 8'd87; b = 8'd178;  #10 
a = 8'd87; b = 8'd179;  #10 
a = 8'd87; b = 8'd180;  #10 
a = 8'd87; b = 8'd181;  #10 
a = 8'd87; b = 8'd182;  #10 
a = 8'd87; b = 8'd183;  #10 
a = 8'd87; b = 8'd184;  #10 
a = 8'd87; b = 8'd185;  #10 
a = 8'd87; b = 8'd186;  #10 
a = 8'd87; b = 8'd187;  #10 
a = 8'd87; b = 8'd188;  #10 
a = 8'd87; b = 8'd189;  #10 
a = 8'd87; b = 8'd190;  #10 
a = 8'd87; b = 8'd191;  #10 
a = 8'd87; b = 8'd192;  #10 
a = 8'd87; b = 8'd193;  #10 
a = 8'd87; b = 8'd194;  #10 
a = 8'd87; b = 8'd195;  #10 
a = 8'd87; b = 8'd196;  #10 
a = 8'd87; b = 8'd197;  #10 
a = 8'd87; b = 8'd198;  #10 
a = 8'd87; b = 8'd199;  #10 
a = 8'd87; b = 8'd200;  #10 
a = 8'd87; b = 8'd201;  #10 
a = 8'd87; b = 8'd202;  #10 
a = 8'd87; b = 8'd203;  #10 
a = 8'd87; b = 8'd204;  #10 
a = 8'd87; b = 8'd205;  #10 
a = 8'd87; b = 8'd206;  #10 
a = 8'd87; b = 8'd207;  #10 
a = 8'd87; b = 8'd208;  #10 
a = 8'd87; b = 8'd209;  #10 
a = 8'd87; b = 8'd210;  #10 
a = 8'd87; b = 8'd211;  #10 
a = 8'd87; b = 8'd212;  #10 
a = 8'd87; b = 8'd213;  #10 
a = 8'd87; b = 8'd214;  #10 
a = 8'd87; b = 8'd215;  #10 
a = 8'd87; b = 8'd216;  #10 
a = 8'd87; b = 8'd217;  #10 
a = 8'd87; b = 8'd218;  #10 
a = 8'd87; b = 8'd219;  #10 
a = 8'd87; b = 8'd220;  #10 
a = 8'd87; b = 8'd221;  #10 
a = 8'd87; b = 8'd222;  #10 
a = 8'd87; b = 8'd223;  #10 
a = 8'd87; b = 8'd224;  #10 
a = 8'd87; b = 8'd225;  #10 
a = 8'd87; b = 8'd226;  #10 
a = 8'd87; b = 8'd227;  #10 
a = 8'd87; b = 8'd228;  #10 
a = 8'd87; b = 8'd229;  #10 
a = 8'd87; b = 8'd230;  #10 
a = 8'd87; b = 8'd231;  #10 
a = 8'd87; b = 8'd232;  #10 
a = 8'd87; b = 8'd233;  #10 
a = 8'd87; b = 8'd234;  #10 
a = 8'd87; b = 8'd235;  #10 
a = 8'd87; b = 8'd236;  #10 
a = 8'd87; b = 8'd237;  #10 
a = 8'd87; b = 8'd238;  #10 
a = 8'd87; b = 8'd239;  #10 
a = 8'd87; b = 8'd240;  #10 
a = 8'd87; b = 8'd241;  #10 
a = 8'd87; b = 8'd242;  #10 
a = 8'd87; b = 8'd243;  #10 
a = 8'd87; b = 8'd244;  #10 
a = 8'd87; b = 8'd245;  #10 
a = 8'd87; b = 8'd246;  #10 
a = 8'd87; b = 8'd247;  #10 
a = 8'd87; b = 8'd248;  #10 
a = 8'd87; b = 8'd249;  #10 
a = 8'd87; b = 8'd250;  #10 
a = 8'd87; b = 8'd251;  #10 
a = 8'd87; b = 8'd252;  #10 
a = 8'd87; b = 8'd253;  #10 
a = 8'd87; b = 8'd254;  #10 
a = 8'd87; b = 8'd255;  #10 
a = 8'd88; b = 8'd0;  #10 
a = 8'd88; b = 8'd1;  #10 
a = 8'd88; b = 8'd2;  #10 
a = 8'd88; b = 8'd3;  #10 
a = 8'd88; b = 8'd4;  #10 
a = 8'd88; b = 8'd5;  #10 
a = 8'd88; b = 8'd6;  #10 
a = 8'd88; b = 8'd7;  #10 
a = 8'd88; b = 8'd8;  #10 
a = 8'd88; b = 8'd9;  #10 
a = 8'd88; b = 8'd10;  #10 
a = 8'd88; b = 8'd11;  #10 
a = 8'd88; b = 8'd12;  #10 
a = 8'd88; b = 8'd13;  #10 
a = 8'd88; b = 8'd14;  #10 
a = 8'd88; b = 8'd15;  #10 
a = 8'd88; b = 8'd16;  #10 
a = 8'd88; b = 8'd17;  #10 
a = 8'd88; b = 8'd18;  #10 
a = 8'd88; b = 8'd19;  #10 
a = 8'd88; b = 8'd20;  #10 
a = 8'd88; b = 8'd21;  #10 
a = 8'd88; b = 8'd22;  #10 
a = 8'd88; b = 8'd23;  #10 
a = 8'd88; b = 8'd24;  #10 
a = 8'd88; b = 8'd25;  #10 
a = 8'd88; b = 8'd26;  #10 
a = 8'd88; b = 8'd27;  #10 
a = 8'd88; b = 8'd28;  #10 
a = 8'd88; b = 8'd29;  #10 
a = 8'd88; b = 8'd30;  #10 
a = 8'd88; b = 8'd31;  #10 
a = 8'd88; b = 8'd32;  #10 
a = 8'd88; b = 8'd33;  #10 
a = 8'd88; b = 8'd34;  #10 
a = 8'd88; b = 8'd35;  #10 
a = 8'd88; b = 8'd36;  #10 
a = 8'd88; b = 8'd37;  #10 
a = 8'd88; b = 8'd38;  #10 
a = 8'd88; b = 8'd39;  #10 
a = 8'd88; b = 8'd40;  #10 
a = 8'd88; b = 8'd41;  #10 
a = 8'd88; b = 8'd42;  #10 
a = 8'd88; b = 8'd43;  #10 
a = 8'd88; b = 8'd44;  #10 
a = 8'd88; b = 8'd45;  #10 
a = 8'd88; b = 8'd46;  #10 
a = 8'd88; b = 8'd47;  #10 
a = 8'd88; b = 8'd48;  #10 
a = 8'd88; b = 8'd49;  #10 
a = 8'd88; b = 8'd50;  #10 
a = 8'd88; b = 8'd51;  #10 
a = 8'd88; b = 8'd52;  #10 
a = 8'd88; b = 8'd53;  #10 
a = 8'd88; b = 8'd54;  #10 
a = 8'd88; b = 8'd55;  #10 
a = 8'd88; b = 8'd56;  #10 
a = 8'd88; b = 8'd57;  #10 
a = 8'd88; b = 8'd58;  #10 
a = 8'd88; b = 8'd59;  #10 
a = 8'd88; b = 8'd60;  #10 
a = 8'd88; b = 8'd61;  #10 
a = 8'd88; b = 8'd62;  #10 
a = 8'd88; b = 8'd63;  #10 
a = 8'd88; b = 8'd64;  #10 
a = 8'd88; b = 8'd65;  #10 
a = 8'd88; b = 8'd66;  #10 
a = 8'd88; b = 8'd67;  #10 
a = 8'd88; b = 8'd68;  #10 
a = 8'd88; b = 8'd69;  #10 
a = 8'd88; b = 8'd70;  #10 
a = 8'd88; b = 8'd71;  #10 
a = 8'd88; b = 8'd72;  #10 
a = 8'd88; b = 8'd73;  #10 
a = 8'd88; b = 8'd74;  #10 
a = 8'd88; b = 8'd75;  #10 
a = 8'd88; b = 8'd76;  #10 
a = 8'd88; b = 8'd77;  #10 
a = 8'd88; b = 8'd78;  #10 
a = 8'd88; b = 8'd79;  #10 
a = 8'd88; b = 8'd80;  #10 
a = 8'd88; b = 8'd81;  #10 
a = 8'd88; b = 8'd82;  #10 
a = 8'd88; b = 8'd83;  #10 
a = 8'd88; b = 8'd84;  #10 
a = 8'd88; b = 8'd85;  #10 
a = 8'd88; b = 8'd86;  #10 
a = 8'd88; b = 8'd87;  #10 
a = 8'd88; b = 8'd88;  #10 
a = 8'd88; b = 8'd89;  #10 
a = 8'd88; b = 8'd90;  #10 
a = 8'd88; b = 8'd91;  #10 
a = 8'd88; b = 8'd92;  #10 
a = 8'd88; b = 8'd93;  #10 
a = 8'd88; b = 8'd94;  #10 
a = 8'd88; b = 8'd95;  #10 
a = 8'd88; b = 8'd96;  #10 
a = 8'd88; b = 8'd97;  #10 
a = 8'd88; b = 8'd98;  #10 
a = 8'd88; b = 8'd99;  #10 
a = 8'd88; b = 8'd100;  #10 
a = 8'd88; b = 8'd101;  #10 
a = 8'd88; b = 8'd102;  #10 
a = 8'd88; b = 8'd103;  #10 
a = 8'd88; b = 8'd104;  #10 
a = 8'd88; b = 8'd105;  #10 
a = 8'd88; b = 8'd106;  #10 
a = 8'd88; b = 8'd107;  #10 
a = 8'd88; b = 8'd108;  #10 
a = 8'd88; b = 8'd109;  #10 
a = 8'd88; b = 8'd110;  #10 
a = 8'd88; b = 8'd111;  #10 
a = 8'd88; b = 8'd112;  #10 
a = 8'd88; b = 8'd113;  #10 
a = 8'd88; b = 8'd114;  #10 
a = 8'd88; b = 8'd115;  #10 
a = 8'd88; b = 8'd116;  #10 
a = 8'd88; b = 8'd117;  #10 
a = 8'd88; b = 8'd118;  #10 
a = 8'd88; b = 8'd119;  #10 
a = 8'd88; b = 8'd120;  #10 
a = 8'd88; b = 8'd121;  #10 
a = 8'd88; b = 8'd122;  #10 
a = 8'd88; b = 8'd123;  #10 
a = 8'd88; b = 8'd124;  #10 
a = 8'd88; b = 8'd125;  #10 
a = 8'd88; b = 8'd126;  #10 
a = 8'd88; b = 8'd127;  #10 
a = 8'd88; b = 8'd128;  #10 
a = 8'd88; b = 8'd129;  #10 
a = 8'd88; b = 8'd130;  #10 
a = 8'd88; b = 8'd131;  #10 
a = 8'd88; b = 8'd132;  #10 
a = 8'd88; b = 8'd133;  #10 
a = 8'd88; b = 8'd134;  #10 
a = 8'd88; b = 8'd135;  #10 
a = 8'd88; b = 8'd136;  #10 
a = 8'd88; b = 8'd137;  #10 
a = 8'd88; b = 8'd138;  #10 
a = 8'd88; b = 8'd139;  #10 
a = 8'd88; b = 8'd140;  #10 
a = 8'd88; b = 8'd141;  #10 
a = 8'd88; b = 8'd142;  #10 
a = 8'd88; b = 8'd143;  #10 
a = 8'd88; b = 8'd144;  #10 
a = 8'd88; b = 8'd145;  #10 
a = 8'd88; b = 8'd146;  #10 
a = 8'd88; b = 8'd147;  #10 
a = 8'd88; b = 8'd148;  #10 
a = 8'd88; b = 8'd149;  #10 
a = 8'd88; b = 8'd150;  #10 
a = 8'd88; b = 8'd151;  #10 
a = 8'd88; b = 8'd152;  #10 
a = 8'd88; b = 8'd153;  #10 
a = 8'd88; b = 8'd154;  #10 
a = 8'd88; b = 8'd155;  #10 
a = 8'd88; b = 8'd156;  #10 
a = 8'd88; b = 8'd157;  #10 
a = 8'd88; b = 8'd158;  #10 
a = 8'd88; b = 8'd159;  #10 
a = 8'd88; b = 8'd160;  #10 
a = 8'd88; b = 8'd161;  #10 
a = 8'd88; b = 8'd162;  #10 
a = 8'd88; b = 8'd163;  #10 
a = 8'd88; b = 8'd164;  #10 
a = 8'd88; b = 8'd165;  #10 
a = 8'd88; b = 8'd166;  #10 
a = 8'd88; b = 8'd167;  #10 
a = 8'd88; b = 8'd168;  #10 
a = 8'd88; b = 8'd169;  #10 
a = 8'd88; b = 8'd170;  #10 
a = 8'd88; b = 8'd171;  #10 
a = 8'd88; b = 8'd172;  #10 
a = 8'd88; b = 8'd173;  #10 
a = 8'd88; b = 8'd174;  #10 
a = 8'd88; b = 8'd175;  #10 
a = 8'd88; b = 8'd176;  #10 
a = 8'd88; b = 8'd177;  #10 
a = 8'd88; b = 8'd178;  #10 
a = 8'd88; b = 8'd179;  #10 
a = 8'd88; b = 8'd180;  #10 
a = 8'd88; b = 8'd181;  #10 
a = 8'd88; b = 8'd182;  #10 
a = 8'd88; b = 8'd183;  #10 
a = 8'd88; b = 8'd184;  #10 
a = 8'd88; b = 8'd185;  #10 
a = 8'd88; b = 8'd186;  #10 
a = 8'd88; b = 8'd187;  #10 
a = 8'd88; b = 8'd188;  #10 
a = 8'd88; b = 8'd189;  #10 
a = 8'd88; b = 8'd190;  #10 
a = 8'd88; b = 8'd191;  #10 
a = 8'd88; b = 8'd192;  #10 
a = 8'd88; b = 8'd193;  #10 
a = 8'd88; b = 8'd194;  #10 
a = 8'd88; b = 8'd195;  #10 
a = 8'd88; b = 8'd196;  #10 
a = 8'd88; b = 8'd197;  #10 
a = 8'd88; b = 8'd198;  #10 
a = 8'd88; b = 8'd199;  #10 
a = 8'd88; b = 8'd200;  #10 
a = 8'd88; b = 8'd201;  #10 
a = 8'd88; b = 8'd202;  #10 
a = 8'd88; b = 8'd203;  #10 
a = 8'd88; b = 8'd204;  #10 
a = 8'd88; b = 8'd205;  #10 
a = 8'd88; b = 8'd206;  #10 
a = 8'd88; b = 8'd207;  #10 
a = 8'd88; b = 8'd208;  #10 
a = 8'd88; b = 8'd209;  #10 
a = 8'd88; b = 8'd210;  #10 
a = 8'd88; b = 8'd211;  #10 
a = 8'd88; b = 8'd212;  #10 
a = 8'd88; b = 8'd213;  #10 
a = 8'd88; b = 8'd214;  #10 
a = 8'd88; b = 8'd215;  #10 
a = 8'd88; b = 8'd216;  #10 
a = 8'd88; b = 8'd217;  #10 
a = 8'd88; b = 8'd218;  #10 
a = 8'd88; b = 8'd219;  #10 
a = 8'd88; b = 8'd220;  #10 
a = 8'd88; b = 8'd221;  #10 
a = 8'd88; b = 8'd222;  #10 
a = 8'd88; b = 8'd223;  #10 
a = 8'd88; b = 8'd224;  #10 
a = 8'd88; b = 8'd225;  #10 
a = 8'd88; b = 8'd226;  #10 
a = 8'd88; b = 8'd227;  #10 
a = 8'd88; b = 8'd228;  #10 
a = 8'd88; b = 8'd229;  #10 
a = 8'd88; b = 8'd230;  #10 
a = 8'd88; b = 8'd231;  #10 
a = 8'd88; b = 8'd232;  #10 
a = 8'd88; b = 8'd233;  #10 
a = 8'd88; b = 8'd234;  #10 
a = 8'd88; b = 8'd235;  #10 
a = 8'd88; b = 8'd236;  #10 
a = 8'd88; b = 8'd237;  #10 
a = 8'd88; b = 8'd238;  #10 
a = 8'd88; b = 8'd239;  #10 
a = 8'd88; b = 8'd240;  #10 
a = 8'd88; b = 8'd241;  #10 
a = 8'd88; b = 8'd242;  #10 
a = 8'd88; b = 8'd243;  #10 
a = 8'd88; b = 8'd244;  #10 
a = 8'd88; b = 8'd245;  #10 
a = 8'd88; b = 8'd246;  #10 
a = 8'd88; b = 8'd247;  #10 
a = 8'd88; b = 8'd248;  #10 
a = 8'd88; b = 8'd249;  #10 
a = 8'd88; b = 8'd250;  #10 
a = 8'd88; b = 8'd251;  #10 
a = 8'd88; b = 8'd252;  #10 
a = 8'd88; b = 8'd253;  #10 
a = 8'd88; b = 8'd254;  #10 
a = 8'd88; b = 8'd255;  #10 
a = 8'd89; b = 8'd0;  #10 
a = 8'd89; b = 8'd1;  #10 
a = 8'd89; b = 8'd2;  #10 
a = 8'd89; b = 8'd3;  #10 
a = 8'd89; b = 8'd4;  #10 
a = 8'd89; b = 8'd5;  #10 
a = 8'd89; b = 8'd6;  #10 
a = 8'd89; b = 8'd7;  #10 
a = 8'd89; b = 8'd8;  #10 
a = 8'd89; b = 8'd9;  #10 
a = 8'd89; b = 8'd10;  #10 
a = 8'd89; b = 8'd11;  #10 
a = 8'd89; b = 8'd12;  #10 
a = 8'd89; b = 8'd13;  #10 
a = 8'd89; b = 8'd14;  #10 
a = 8'd89; b = 8'd15;  #10 
a = 8'd89; b = 8'd16;  #10 
a = 8'd89; b = 8'd17;  #10 
a = 8'd89; b = 8'd18;  #10 
a = 8'd89; b = 8'd19;  #10 
a = 8'd89; b = 8'd20;  #10 
a = 8'd89; b = 8'd21;  #10 
a = 8'd89; b = 8'd22;  #10 
a = 8'd89; b = 8'd23;  #10 
a = 8'd89; b = 8'd24;  #10 
a = 8'd89; b = 8'd25;  #10 
a = 8'd89; b = 8'd26;  #10 
a = 8'd89; b = 8'd27;  #10 
a = 8'd89; b = 8'd28;  #10 
a = 8'd89; b = 8'd29;  #10 
a = 8'd89; b = 8'd30;  #10 
a = 8'd89; b = 8'd31;  #10 
a = 8'd89; b = 8'd32;  #10 
a = 8'd89; b = 8'd33;  #10 
a = 8'd89; b = 8'd34;  #10 
a = 8'd89; b = 8'd35;  #10 
a = 8'd89; b = 8'd36;  #10 
a = 8'd89; b = 8'd37;  #10 
a = 8'd89; b = 8'd38;  #10 
a = 8'd89; b = 8'd39;  #10 
a = 8'd89; b = 8'd40;  #10 
a = 8'd89; b = 8'd41;  #10 
a = 8'd89; b = 8'd42;  #10 
a = 8'd89; b = 8'd43;  #10 
a = 8'd89; b = 8'd44;  #10 
a = 8'd89; b = 8'd45;  #10 
a = 8'd89; b = 8'd46;  #10 
a = 8'd89; b = 8'd47;  #10 
a = 8'd89; b = 8'd48;  #10 
a = 8'd89; b = 8'd49;  #10 
a = 8'd89; b = 8'd50;  #10 
a = 8'd89; b = 8'd51;  #10 
a = 8'd89; b = 8'd52;  #10 
a = 8'd89; b = 8'd53;  #10 
a = 8'd89; b = 8'd54;  #10 
a = 8'd89; b = 8'd55;  #10 
a = 8'd89; b = 8'd56;  #10 
a = 8'd89; b = 8'd57;  #10 
a = 8'd89; b = 8'd58;  #10 
a = 8'd89; b = 8'd59;  #10 
a = 8'd89; b = 8'd60;  #10 
a = 8'd89; b = 8'd61;  #10 
a = 8'd89; b = 8'd62;  #10 
a = 8'd89; b = 8'd63;  #10 
a = 8'd89; b = 8'd64;  #10 
a = 8'd89; b = 8'd65;  #10 
a = 8'd89; b = 8'd66;  #10 
a = 8'd89; b = 8'd67;  #10 
a = 8'd89; b = 8'd68;  #10 
a = 8'd89; b = 8'd69;  #10 
a = 8'd89; b = 8'd70;  #10 
a = 8'd89; b = 8'd71;  #10 
a = 8'd89; b = 8'd72;  #10 
a = 8'd89; b = 8'd73;  #10 
a = 8'd89; b = 8'd74;  #10 
a = 8'd89; b = 8'd75;  #10 
a = 8'd89; b = 8'd76;  #10 
a = 8'd89; b = 8'd77;  #10 
a = 8'd89; b = 8'd78;  #10 
a = 8'd89; b = 8'd79;  #10 
a = 8'd89; b = 8'd80;  #10 
a = 8'd89; b = 8'd81;  #10 
a = 8'd89; b = 8'd82;  #10 
a = 8'd89; b = 8'd83;  #10 
a = 8'd89; b = 8'd84;  #10 
a = 8'd89; b = 8'd85;  #10 
a = 8'd89; b = 8'd86;  #10 
a = 8'd89; b = 8'd87;  #10 
a = 8'd89; b = 8'd88;  #10 
a = 8'd89; b = 8'd89;  #10 
a = 8'd89; b = 8'd90;  #10 
a = 8'd89; b = 8'd91;  #10 
a = 8'd89; b = 8'd92;  #10 
a = 8'd89; b = 8'd93;  #10 
a = 8'd89; b = 8'd94;  #10 
a = 8'd89; b = 8'd95;  #10 
a = 8'd89; b = 8'd96;  #10 
a = 8'd89; b = 8'd97;  #10 
a = 8'd89; b = 8'd98;  #10 
a = 8'd89; b = 8'd99;  #10 
a = 8'd89; b = 8'd100;  #10 
a = 8'd89; b = 8'd101;  #10 
a = 8'd89; b = 8'd102;  #10 
a = 8'd89; b = 8'd103;  #10 
a = 8'd89; b = 8'd104;  #10 
a = 8'd89; b = 8'd105;  #10 
a = 8'd89; b = 8'd106;  #10 
a = 8'd89; b = 8'd107;  #10 
a = 8'd89; b = 8'd108;  #10 
a = 8'd89; b = 8'd109;  #10 
a = 8'd89; b = 8'd110;  #10 
a = 8'd89; b = 8'd111;  #10 
a = 8'd89; b = 8'd112;  #10 
a = 8'd89; b = 8'd113;  #10 
a = 8'd89; b = 8'd114;  #10 
a = 8'd89; b = 8'd115;  #10 
a = 8'd89; b = 8'd116;  #10 
a = 8'd89; b = 8'd117;  #10 
a = 8'd89; b = 8'd118;  #10 
a = 8'd89; b = 8'd119;  #10 
a = 8'd89; b = 8'd120;  #10 
a = 8'd89; b = 8'd121;  #10 
a = 8'd89; b = 8'd122;  #10 
a = 8'd89; b = 8'd123;  #10 
a = 8'd89; b = 8'd124;  #10 
a = 8'd89; b = 8'd125;  #10 
a = 8'd89; b = 8'd126;  #10 
a = 8'd89; b = 8'd127;  #10 
a = 8'd89; b = 8'd128;  #10 
a = 8'd89; b = 8'd129;  #10 
a = 8'd89; b = 8'd130;  #10 
a = 8'd89; b = 8'd131;  #10 
a = 8'd89; b = 8'd132;  #10 
a = 8'd89; b = 8'd133;  #10 
a = 8'd89; b = 8'd134;  #10 
a = 8'd89; b = 8'd135;  #10 
a = 8'd89; b = 8'd136;  #10 
a = 8'd89; b = 8'd137;  #10 
a = 8'd89; b = 8'd138;  #10 
a = 8'd89; b = 8'd139;  #10 
a = 8'd89; b = 8'd140;  #10 
a = 8'd89; b = 8'd141;  #10 
a = 8'd89; b = 8'd142;  #10 
a = 8'd89; b = 8'd143;  #10 
a = 8'd89; b = 8'd144;  #10 
a = 8'd89; b = 8'd145;  #10 
a = 8'd89; b = 8'd146;  #10 
a = 8'd89; b = 8'd147;  #10 
a = 8'd89; b = 8'd148;  #10 
a = 8'd89; b = 8'd149;  #10 
a = 8'd89; b = 8'd150;  #10 
a = 8'd89; b = 8'd151;  #10 
a = 8'd89; b = 8'd152;  #10 
a = 8'd89; b = 8'd153;  #10 
a = 8'd89; b = 8'd154;  #10 
a = 8'd89; b = 8'd155;  #10 
a = 8'd89; b = 8'd156;  #10 
a = 8'd89; b = 8'd157;  #10 
a = 8'd89; b = 8'd158;  #10 
a = 8'd89; b = 8'd159;  #10 
a = 8'd89; b = 8'd160;  #10 
a = 8'd89; b = 8'd161;  #10 
a = 8'd89; b = 8'd162;  #10 
a = 8'd89; b = 8'd163;  #10 
a = 8'd89; b = 8'd164;  #10 
a = 8'd89; b = 8'd165;  #10 
a = 8'd89; b = 8'd166;  #10 
a = 8'd89; b = 8'd167;  #10 
a = 8'd89; b = 8'd168;  #10 
a = 8'd89; b = 8'd169;  #10 
a = 8'd89; b = 8'd170;  #10 
a = 8'd89; b = 8'd171;  #10 
a = 8'd89; b = 8'd172;  #10 
a = 8'd89; b = 8'd173;  #10 
a = 8'd89; b = 8'd174;  #10 
a = 8'd89; b = 8'd175;  #10 
a = 8'd89; b = 8'd176;  #10 
a = 8'd89; b = 8'd177;  #10 
a = 8'd89; b = 8'd178;  #10 
a = 8'd89; b = 8'd179;  #10 
a = 8'd89; b = 8'd180;  #10 
a = 8'd89; b = 8'd181;  #10 
a = 8'd89; b = 8'd182;  #10 
a = 8'd89; b = 8'd183;  #10 
a = 8'd89; b = 8'd184;  #10 
a = 8'd89; b = 8'd185;  #10 
a = 8'd89; b = 8'd186;  #10 
a = 8'd89; b = 8'd187;  #10 
a = 8'd89; b = 8'd188;  #10 
a = 8'd89; b = 8'd189;  #10 
a = 8'd89; b = 8'd190;  #10 
a = 8'd89; b = 8'd191;  #10 
a = 8'd89; b = 8'd192;  #10 
a = 8'd89; b = 8'd193;  #10 
a = 8'd89; b = 8'd194;  #10 
a = 8'd89; b = 8'd195;  #10 
a = 8'd89; b = 8'd196;  #10 
a = 8'd89; b = 8'd197;  #10 
a = 8'd89; b = 8'd198;  #10 
a = 8'd89; b = 8'd199;  #10 
a = 8'd89; b = 8'd200;  #10 
a = 8'd89; b = 8'd201;  #10 
a = 8'd89; b = 8'd202;  #10 
a = 8'd89; b = 8'd203;  #10 
a = 8'd89; b = 8'd204;  #10 
a = 8'd89; b = 8'd205;  #10 
a = 8'd89; b = 8'd206;  #10 
a = 8'd89; b = 8'd207;  #10 
a = 8'd89; b = 8'd208;  #10 
a = 8'd89; b = 8'd209;  #10 
a = 8'd89; b = 8'd210;  #10 
a = 8'd89; b = 8'd211;  #10 
a = 8'd89; b = 8'd212;  #10 
a = 8'd89; b = 8'd213;  #10 
a = 8'd89; b = 8'd214;  #10 
a = 8'd89; b = 8'd215;  #10 
a = 8'd89; b = 8'd216;  #10 
a = 8'd89; b = 8'd217;  #10 
a = 8'd89; b = 8'd218;  #10 
a = 8'd89; b = 8'd219;  #10 
a = 8'd89; b = 8'd220;  #10 
a = 8'd89; b = 8'd221;  #10 
a = 8'd89; b = 8'd222;  #10 
a = 8'd89; b = 8'd223;  #10 
a = 8'd89; b = 8'd224;  #10 
a = 8'd89; b = 8'd225;  #10 
a = 8'd89; b = 8'd226;  #10 
a = 8'd89; b = 8'd227;  #10 
a = 8'd89; b = 8'd228;  #10 
a = 8'd89; b = 8'd229;  #10 
a = 8'd89; b = 8'd230;  #10 
a = 8'd89; b = 8'd231;  #10 
a = 8'd89; b = 8'd232;  #10 
a = 8'd89; b = 8'd233;  #10 
a = 8'd89; b = 8'd234;  #10 
a = 8'd89; b = 8'd235;  #10 
a = 8'd89; b = 8'd236;  #10 
a = 8'd89; b = 8'd237;  #10 
a = 8'd89; b = 8'd238;  #10 
a = 8'd89; b = 8'd239;  #10 
a = 8'd89; b = 8'd240;  #10 
a = 8'd89; b = 8'd241;  #10 
a = 8'd89; b = 8'd242;  #10 
a = 8'd89; b = 8'd243;  #10 
a = 8'd89; b = 8'd244;  #10 
a = 8'd89; b = 8'd245;  #10 
a = 8'd89; b = 8'd246;  #10 
a = 8'd89; b = 8'd247;  #10 
a = 8'd89; b = 8'd248;  #10 
a = 8'd89; b = 8'd249;  #10 
a = 8'd89; b = 8'd250;  #10 
a = 8'd89; b = 8'd251;  #10 
a = 8'd89; b = 8'd252;  #10 
a = 8'd89; b = 8'd253;  #10 
a = 8'd89; b = 8'd254;  #10 
a = 8'd89; b = 8'd255;  #10 
a = 8'd90; b = 8'd0;  #10 
a = 8'd90; b = 8'd1;  #10 
a = 8'd90; b = 8'd2;  #10 
a = 8'd90; b = 8'd3;  #10 
a = 8'd90; b = 8'd4;  #10 
a = 8'd90; b = 8'd5;  #10 
a = 8'd90; b = 8'd6;  #10 
a = 8'd90; b = 8'd7;  #10 
a = 8'd90; b = 8'd8;  #10 
a = 8'd90; b = 8'd9;  #10 
a = 8'd90; b = 8'd10;  #10 
a = 8'd90; b = 8'd11;  #10 
a = 8'd90; b = 8'd12;  #10 
a = 8'd90; b = 8'd13;  #10 
a = 8'd90; b = 8'd14;  #10 
a = 8'd90; b = 8'd15;  #10 
a = 8'd90; b = 8'd16;  #10 
a = 8'd90; b = 8'd17;  #10 
a = 8'd90; b = 8'd18;  #10 
a = 8'd90; b = 8'd19;  #10 
a = 8'd90; b = 8'd20;  #10 
a = 8'd90; b = 8'd21;  #10 
a = 8'd90; b = 8'd22;  #10 
a = 8'd90; b = 8'd23;  #10 
a = 8'd90; b = 8'd24;  #10 
a = 8'd90; b = 8'd25;  #10 
a = 8'd90; b = 8'd26;  #10 
a = 8'd90; b = 8'd27;  #10 
a = 8'd90; b = 8'd28;  #10 
a = 8'd90; b = 8'd29;  #10 
a = 8'd90; b = 8'd30;  #10 
a = 8'd90; b = 8'd31;  #10 
a = 8'd90; b = 8'd32;  #10 
a = 8'd90; b = 8'd33;  #10 
a = 8'd90; b = 8'd34;  #10 
a = 8'd90; b = 8'd35;  #10 
a = 8'd90; b = 8'd36;  #10 
a = 8'd90; b = 8'd37;  #10 
a = 8'd90; b = 8'd38;  #10 
a = 8'd90; b = 8'd39;  #10 
a = 8'd90; b = 8'd40;  #10 
a = 8'd90; b = 8'd41;  #10 
a = 8'd90; b = 8'd42;  #10 
a = 8'd90; b = 8'd43;  #10 
a = 8'd90; b = 8'd44;  #10 
a = 8'd90; b = 8'd45;  #10 
a = 8'd90; b = 8'd46;  #10 
a = 8'd90; b = 8'd47;  #10 
a = 8'd90; b = 8'd48;  #10 
a = 8'd90; b = 8'd49;  #10 
a = 8'd90; b = 8'd50;  #10 
a = 8'd90; b = 8'd51;  #10 
a = 8'd90; b = 8'd52;  #10 
a = 8'd90; b = 8'd53;  #10 
a = 8'd90; b = 8'd54;  #10 
a = 8'd90; b = 8'd55;  #10 
a = 8'd90; b = 8'd56;  #10 
a = 8'd90; b = 8'd57;  #10 
a = 8'd90; b = 8'd58;  #10 
a = 8'd90; b = 8'd59;  #10 
a = 8'd90; b = 8'd60;  #10 
a = 8'd90; b = 8'd61;  #10 
a = 8'd90; b = 8'd62;  #10 
a = 8'd90; b = 8'd63;  #10 
a = 8'd90; b = 8'd64;  #10 
a = 8'd90; b = 8'd65;  #10 
a = 8'd90; b = 8'd66;  #10 
a = 8'd90; b = 8'd67;  #10 
a = 8'd90; b = 8'd68;  #10 
a = 8'd90; b = 8'd69;  #10 
a = 8'd90; b = 8'd70;  #10 
a = 8'd90; b = 8'd71;  #10 
a = 8'd90; b = 8'd72;  #10 
a = 8'd90; b = 8'd73;  #10 
a = 8'd90; b = 8'd74;  #10 
a = 8'd90; b = 8'd75;  #10 
a = 8'd90; b = 8'd76;  #10 
a = 8'd90; b = 8'd77;  #10 
a = 8'd90; b = 8'd78;  #10 
a = 8'd90; b = 8'd79;  #10 
a = 8'd90; b = 8'd80;  #10 
a = 8'd90; b = 8'd81;  #10 
a = 8'd90; b = 8'd82;  #10 
a = 8'd90; b = 8'd83;  #10 
a = 8'd90; b = 8'd84;  #10 
a = 8'd90; b = 8'd85;  #10 
a = 8'd90; b = 8'd86;  #10 
a = 8'd90; b = 8'd87;  #10 
a = 8'd90; b = 8'd88;  #10 
a = 8'd90; b = 8'd89;  #10 
a = 8'd90; b = 8'd90;  #10 
a = 8'd90; b = 8'd91;  #10 
a = 8'd90; b = 8'd92;  #10 
a = 8'd90; b = 8'd93;  #10 
a = 8'd90; b = 8'd94;  #10 
a = 8'd90; b = 8'd95;  #10 
a = 8'd90; b = 8'd96;  #10 
a = 8'd90; b = 8'd97;  #10 
a = 8'd90; b = 8'd98;  #10 
a = 8'd90; b = 8'd99;  #10 
a = 8'd90; b = 8'd100;  #10 
a = 8'd90; b = 8'd101;  #10 
a = 8'd90; b = 8'd102;  #10 
a = 8'd90; b = 8'd103;  #10 
a = 8'd90; b = 8'd104;  #10 
a = 8'd90; b = 8'd105;  #10 
a = 8'd90; b = 8'd106;  #10 
a = 8'd90; b = 8'd107;  #10 
a = 8'd90; b = 8'd108;  #10 
a = 8'd90; b = 8'd109;  #10 
a = 8'd90; b = 8'd110;  #10 
a = 8'd90; b = 8'd111;  #10 
a = 8'd90; b = 8'd112;  #10 
a = 8'd90; b = 8'd113;  #10 
a = 8'd90; b = 8'd114;  #10 
a = 8'd90; b = 8'd115;  #10 
a = 8'd90; b = 8'd116;  #10 
a = 8'd90; b = 8'd117;  #10 
a = 8'd90; b = 8'd118;  #10 
a = 8'd90; b = 8'd119;  #10 
a = 8'd90; b = 8'd120;  #10 
a = 8'd90; b = 8'd121;  #10 
a = 8'd90; b = 8'd122;  #10 
a = 8'd90; b = 8'd123;  #10 
a = 8'd90; b = 8'd124;  #10 
a = 8'd90; b = 8'd125;  #10 
a = 8'd90; b = 8'd126;  #10 
a = 8'd90; b = 8'd127;  #10 
a = 8'd90; b = 8'd128;  #10 
a = 8'd90; b = 8'd129;  #10 
a = 8'd90; b = 8'd130;  #10 
a = 8'd90; b = 8'd131;  #10 
a = 8'd90; b = 8'd132;  #10 
a = 8'd90; b = 8'd133;  #10 
a = 8'd90; b = 8'd134;  #10 
a = 8'd90; b = 8'd135;  #10 
a = 8'd90; b = 8'd136;  #10 
a = 8'd90; b = 8'd137;  #10 
a = 8'd90; b = 8'd138;  #10 
a = 8'd90; b = 8'd139;  #10 
a = 8'd90; b = 8'd140;  #10 
a = 8'd90; b = 8'd141;  #10 
a = 8'd90; b = 8'd142;  #10 
a = 8'd90; b = 8'd143;  #10 
a = 8'd90; b = 8'd144;  #10 
a = 8'd90; b = 8'd145;  #10 
a = 8'd90; b = 8'd146;  #10 
a = 8'd90; b = 8'd147;  #10 
a = 8'd90; b = 8'd148;  #10 
a = 8'd90; b = 8'd149;  #10 
a = 8'd90; b = 8'd150;  #10 
a = 8'd90; b = 8'd151;  #10 
a = 8'd90; b = 8'd152;  #10 
a = 8'd90; b = 8'd153;  #10 
a = 8'd90; b = 8'd154;  #10 
a = 8'd90; b = 8'd155;  #10 
a = 8'd90; b = 8'd156;  #10 
a = 8'd90; b = 8'd157;  #10 
a = 8'd90; b = 8'd158;  #10 
a = 8'd90; b = 8'd159;  #10 
a = 8'd90; b = 8'd160;  #10 
a = 8'd90; b = 8'd161;  #10 
a = 8'd90; b = 8'd162;  #10 
a = 8'd90; b = 8'd163;  #10 
a = 8'd90; b = 8'd164;  #10 
a = 8'd90; b = 8'd165;  #10 
a = 8'd90; b = 8'd166;  #10 
a = 8'd90; b = 8'd167;  #10 
a = 8'd90; b = 8'd168;  #10 
a = 8'd90; b = 8'd169;  #10 
a = 8'd90; b = 8'd170;  #10 
a = 8'd90; b = 8'd171;  #10 
a = 8'd90; b = 8'd172;  #10 
a = 8'd90; b = 8'd173;  #10 
a = 8'd90; b = 8'd174;  #10 
a = 8'd90; b = 8'd175;  #10 
a = 8'd90; b = 8'd176;  #10 
a = 8'd90; b = 8'd177;  #10 
a = 8'd90; b = 8'd178;  #10 
a = 8'd90; b = 8'd179;  #10 
a = 8'd90; b = 8'd180;  #10 
a = 8'd90; b = 8'd181;  #10 
a = 8'd90; b = 8'd182;  #10 
a = 8'd90; b = 8'd183;  #10 
a = 8'd90; b = 8'd184;  #10 
a = 8'd90; b = 8'd185;  #10 
a = 8'd90; b = 8'd186;  #10 
a = 8'd90; b = 8'd187;  #10 
a = 8'd90; b = 8'd188;  #10 
a = 8'd90; b = 8'd189;  #10 
a = 8'd90; b = 8'd190;  #10 
a = 8'd90; b = 8'd191;  #10 
a = 8'd90; b = 8'd192;  #10 
a = 8'd90; b = 8'd193;  #10 
a = 8'd90; b = 8'd194;  #10 
a = 8'd90; b = 8'd195;  #10 
a = 8'd90; b = 8'd196;  #10 
a = 8'd90; b = 8'd197;  #10 
a = 8'd90; b = 8'd198;  #10 
a = 8'd90; b = 8'd199;  #10 
a = 8'd90; b = 8'd200;  #10 
a = 8'd90; b = 8'd201;  #10 
a = 8'd90; b = 8'd202;  #10 
a = 8'd90; b = 8'd203;  #10 
a = 8'd90; b = 8'd204;  #10 
a = 8'd90; b = 8'd205;  #10 
a = 8'd90; b = 8'd206;  #10 
a = 8'd90; b = 8'd207;  #10 
a = 8'd90; b = 8'd208;  #10 
a = 8'd90; b = 8'd209;  #10 
a = 8'd90; b = 8'd210;  #10 
a = 8'd90; b = 8'd211;  #10 
a = 8'd90; b = 8'd212;  #10 
a = 8'd90; b = 8'd213;  #10 
a = 8'd90; b = 8'd214;  #10 
a = 8'd90; b = 8'd215;  #10 
a = 8'd90; b = 8'd216;  #10 
a = 8'd90; b = 8'd217;  #10 
a = 8'd90; b = 8'd218;  #10 
a = 8'd90; b = 8'd219;  #10 
a = 8'd90; b = 8'd220;  #10 
a = 8'd90; b = 8'd221;  #10 
a = 8'd90; b = 8'd222;  #10 
a = 8'd90; b = 8'd223;  #10 
a = 8'd90; b = 8'd224;  #10 
a = 8'd90; b = 8'd225;  #10 
a = 8'd90; b = 8'd226;  #10 
a = 8'd90; b = 8'd227;  #10 
a = 8'd90; b = 8'd228;  #10 
a = 8'd90; b = 8'd229;  #10 
a = 8'd90; b = 8'd230;  #10 
a = 8'd90; b = 8'd231;  #10 
a = 8'd90; b = 8'd232;  #10 
a = 8'd90; b = 8'd233;  #10 
a = 8'd90; b = 8'd234;  #10 
a = 8'd90; b = 8'd235;  #10 
a = 8'd90; b = 8'd236;  #10 
a = 8'd90; b = 8'd237;  #10 
a = 8'd90; b = 8'd238;  #10 
a = 8'd90; b = 8'd239;  #10 
a = 8'd90; b = 8'd240;  #10 
a = 8'd90; b = 8'd241;  #10 
a = 8'd90; b = 8'd242;  #10 
a = 8'd90; b = 8'd243;  #10 
a = 8'd90; b = 8'd244;  #10 
a = 8'd90; b = 8'd245;  #10 
a = 8'd90; b = 8'd246;  #10 
a = 8'd90; b = 8'd247;  #10 
a = 8'd90; b = 8'd248;  #10 
a = 8'd90; b = 8'd249;  #10 
a = 8'd90; b = 8'd250;  #10 
a = 8'd90; b = 8'd251;  #10 
a = 8'd90; b = 8'd252;  #10 
a = 8'd90; b = 8'd253;  #10 
a = 8'd90; b = 8'd254;  #10 
a = 8'd90; b = 8'd255;  #10 
a = 8'd91; b = 8'd0;  #10 
a = 8'd91; b = 8'd1;  #10 
a = 8'd91; b = 8'd2;  #10 
a = 8'd91; b = 8'd3;  #10 
a = 8'd91; b = 8'd4;  #10 
a = 8'd91; b = 8'd5;  #10 
a = 8'd91; b = 8'd6;  #10 
a = 8'd91; b = 8'd7;  #10 
a = 8'd91; b = 8'd8;  #10 
a = 8'd91; b = 8'd9;  #10 
a = 8'd91; b = 8'd10;  #10 
a = 8'd91; b = 8'd11;  #10 
a = 8'd91; b = 8'd12;  #10 
a = 8'd91; b = 8'd13;  #10 
a = 8'd91; b = 8'd14;  #10 
a = 8'd91; b = 8'd15;  #10 
a = 8'd91; b = 8'd16;  #10 
a = 8'd91; b = 8'd17;  #10 
a = 8'd91; b = 8'd18;  #10 
a = 8'd91; b = 8'd19;  #10 
a = 8'd91; b = 8'd20;  #10 
a = 8'd91; b = 8'd21;  #10 
a = 8'd91; b = 8'd22;  #10 
a = 8'd91; b = 8'd23;  #10 
a = 8'd91; b = 8'd24;  #10 
a = 8'd91; b = 8'd25;  #10 
a = 8'd91; b = 8'd26;  #10 
a = 8'd91; b = 8'd27;  #10 
a = 8'd91; b = 8'd28;  #10 
a = 8'd91; b = 8'd29;  #10 
a = 8'd91; b = 8'd30;  #10 
a = 8'd91; b = 8'd31;  #10 
a = 8'd91; b = 8'd32;  #10 
a = 8'd91; b = 8'd33;  #10 
a = 8'd91; b = 8'd34;  #10 
a = 8'd91; b = 8'd35;  #10 
a = 8'd91; b = 8'd36;  #10 
a = 8'd91; b = 8'd37;  #10 
a = 8'd91; b = 8'd38;  #10 
a = 8'd91; b = 8'd39;  #10 
a = 8'd91; b = 8'd40;  #10 
a = 8'd91; b = 8'd41;  #10 
a = 8'd91; b = 8'd42;  #10 
a = 8'd91; b = 8'd43;  #10 
a = 8'd91; b = 8'd44;  #10 
a = 8'd91; b = 8'd45;  #10 
a = 8'd91; b = 8'd46;  #10 
a = 8'd91; b = 8'd47;  #10 
a = 8'd91; b = 8'd48;  #10 
a = 8'd91; b = 8'd49;  #10 
a = 8'd91; b = 8'd50;  #10 
a = 8'd91; b = 8'd51;  #10 
a = 8'd91; b = 8'd52;  #10 
a = 8'd91; b = 8'd53;  #10 
a = 8'd91; b = 8'd54;  #10 
a = 8'd91; b = 8'd55;  #10 
a = 8'd91; b = 8'd56;  #10 
a = 8'd91; b = 8'd57;  #10 
a = 8'd91; b = 8'd58;  #10 
a = 8'd91; b = 8'd59;  #10 
a = 8'd91; b = 8'd60;  #10 
a = 8'd91; b = 8'd61;  #10 
a = 8'd91; b = 8'd62;  #10 
a = 8'd91; b = 8'd63;  #10 
a = 8'd91; b = 8'd64;  #10 
a = 8'd91; b = 8'd65;  #10 
a = 8'd91; b = 8'd66;  #10 
a = 8'd91; b = 8'd67;  #10 
a = 8'd91; b = 8'd68;  #10 
a = 8'd91; b = 8'd69;  #10 
a = 8'd91; b = 8'd70;  #10 
a = 8'd91; b = 8'd71;  #10 
a = 8'd91; b = 8'd72;  #10 
a = 8'd91; b = 8'd73;  #10 
a = 8'd91; b = 8'd74;  #10 
a = 8'd91; b = 8'd75;  #10 
a = 8'd91; b = 8'd76;  #10 
a = 8'd91; b = 8'd77;  #10 
a = 8'd91; b = 8'd78;  #10 
a = 8'd91; b = 8'd79;  #10 
a = 8'd91; b = 8'd80;  #10 
a = 8'd91; b = 8'd81;  #10 
a = 8'd91; b = 8'd82;  #10 
a = 8'd91; b = 8'd83;  #10 
a = 8'd91; b = 8'd84;  #10 
a = 8'd91; b = 8'd85;  #10 
a = 8'd91; b = 8'd86;  #10 
a = 8'd91; b = 8'd87;  #10 
a = 8'd91; b = 8'd88;  #10 
a = 8'd91; b = 8'd89;  #10 
a = 8'd91; b = 8'd90;  #10 
a = 8'd91; b = 8'd91;  #10 
a = 8'd91; b = 8'd92;  #10 
a = 8'd91; b = 8'd93;  #10 
a = 8'd91; b = 8'd94;  #10 
a = 8'd91; b = 8'd95;  #10 
a = 8'd91; b = 8'd96;  #10 
a = 8'd91; b = 8'd97;  #10 
a = 8'd91; b = 8'd98;  #10 
a = 8'd91; b = 8'd99;  #10 
a = 8'd91; b = 8'd100;  #10 
a = 8'd91; b = 8'd101;  #10 
a = 8'd91; b = 8'd102;  #10 
a = 8'd91; b = 8'd103;  #10 
a = 8'd91; b = 8'd104;  #10 
a = 8'd91; b = 8'd105;  #10 
a = 8'd91; b = 8'd106;  #10 
a = 8'd91; b = 8'd107;  #10 
a = 8'd91; b = 8'd108;  #10 
a = 8'd91; b = 8'd109;  #10 
a = 8'd91; b = 8'd110;  #10 
a = 8'd91; b = 8'd111;  #10 
a = 8'd91; b = 8'd112;  #10 
a = 8'd91; b = 8'd113;  #10 
a = 8'd91; b = 8'd114;  #10 
a = 8'd91; b = 8'd115;  #10 
a = 8'd91; b = 8'd116;  #10 
a = 8'd91; b = 8'd117;  #10 
a = 8'd91; b = 8'd118;  #10 
a = 8'd91; b = 8'd119;  #10 
a = 8'd91; b = 8'd120;  #10 
a = 8'd91; b = 8'd121;  #10 
a = 8'd91; b = 8'd122;  #10 
a = 8'd91; b = 8'd123;  #10 
a = 8'd91; b = 8'd124;  #10 
a = 8'd91; b = 8'd125;  #10 
a = 8'd91; b = 8'd126;  #10 
a = 8'd91; b = 8'd127;  #10 
a = 8'd91; b = 8'd128;  #10 
a = 8'd91; b = 8'd129;  #10 
a = 8'd91; b = 8'd130;  #10 
a = 8'd91; b = 8'd131;  #10 
a = 8'd91; b = 8'd132;  #10 
a = 8'd91; b = 8'd133;  #10 
a = 8'd91; b = 8'd134;  #10 
a = 8'd91; b = 8'd135;  #10 
a = 8'd91; b = 8'd136;  #10 
a = 8'd91; b = 8'd137;  #10 
a = 8'd91; b = 8'd138;  #10 
a = 8'd91; b = 8'd139;  #10 
a = 8'd91; b = 8'd140;  #10 
a = 8'd91; b = 8'd141;  #10 
a = 8'd91; b = 8'd142;  #10 
a = 8'd91; b = 8'd143;  #10 
a = 8'd91; b = 8'd144;  #10 
a = 8'd91; b = 8'd145;  #10 
a = 8'd91; b = 8'd146;  #10 
a = 8'd91; b = 8'd147;  #10 
a = 8'd91; b = 8'd148;  #10 
a = 8'd91; b = 8'd149;  #10 
a = 8'd91; b = 8'd150;  #10 
a = 8'd91; b = 8'd151;  #10 
a = 8'd91; b = 8'd152;  #10 
a = 8'd91; b = 8'd153;  #10 
a = 8'd91; b = 8'd154;  #10 
a = 8'd91; b = 8'd155;  #10 
a = 8'd91; b = 8'd156;  #10 
a = 8'd91; b = 8'd157;  #10 
a = 8'd91; b = 8'd158;  #10 
a = 8'd91; b = 8'd159;  #10 
a = 8'd91; b = 8'd160;  #10 
a = 8'd91; b = 8'd161;  #10 
a = 8'd91; b = 8'd162;  #10 
a = 8'd91; b = 8'd163;  #10 
a = 8'd91; b = 8'd164;  #10 
a = 8'd91; b = 8'd165;  #10 
a = 8'd91; b = 8'd166;  #10 
a = 8'd91; b = 8'd167;  #10 
a = 8'd91; b = 8'd168;  #10 
a = 8'd91; b = 8'd169;  #10 
a = 8'd91; b = 8'd170;  #10 
a = 8'd91; b = 8'd171;  #10 
a = 8'd91; b = 8'd172;  #10 
a = 8'd91; b = 8'd173;  #10 
a = 8'd91; b = 8'd174;  #10 
a = 8'd91; b = 8'd175;  #10 
a = 8'd91; b = 8'd176;  #10 
a = 8'd91; b = 8'd177;  #10 
a = 8'd91; b = 8'd178;  #10 
a = 8'd91; b = 8'd179;  #10 
a = 8'd91; b = 8'd180;  #10 
a = 8'd91; b = 8'd181;  #10 
a = 8'd91; b = 8'd182;  #10 
a = 8'd91; b = 8'd183;  #10 
a = 8'd91; b = 8'd184;  #10 
a = 8'd91; b = 8'd185;  #10 
a = 8'd91; b = 8'd186;  #10 
a = 8'd91; b = 8'd187;  #10 
a = 8'd91; b = 8'd188;  #10 
a = 8'd91; b = 8'd189;  #10 
a = 8'd91; b = 8'd190;  #10 
a = 8'd91; b = 8'd191;  #10 
a = 8'd91; b = 8'd192;  #10 
a = 8'd91; b = 8'd193;  #10 
a = 8'd91; b = 8'd194;  #10 
a = 8'd91; b = 8'd195;  #10 
a = 8'd91; b = 8'd196;  #10 
a = 8'd91; b = 8'd197;  #10 
a = 8'd91; b = 8'd198;  #10 
a = 8'd91; b = 8'd199;  #10 
a = 8'd91; b = 8'd200;  #10 
a = 8'd91; b = 8'd201;  #10 
a = 8'd91; b = 8'd202;  #10 
a = 8'd91; b = 8'd203;  #10 
a = 8'd91; b = 8'd204;  #10 
a = 8'd91; b = 8'd205;  #10 
a = 8'd91; b = 8'd206;  #10 
a = 8'd91; b = 8'd207;  #10 
a = 8'd91; b = 8'd208;  #10 
a = 8'd91; b = 8'd209;  #10 
a = 8'd91; b = 8'd210;  #10 
a = 8'd91; b = 8'd211;  #10 
a = 8'd91; b = 8'd212;  #10 
a = 8'd91; b = 8'd213;  #10 
a = 8'd91; b = 8'd214;  #10 
a = 8'd91; b = 8'd215;  #10 
a = 8'd91; b = 8'd216;  #10 
a = 8'd91; b = 8'd217;  #10 
a = 8'd91; b = 8'd218;  #10 
a = 8'd91; b = 8'd219;  #10 
a = 8'd91; b = 8'd220;  #10 
a = 8'd91; b = 8'd221;  #10 
a = 8'd91; b = 8'd222;  #10 
a = 8'd91; b = 8'd223;  #10 
a = 8'd91; b = 8'd224;  #10 
a = 8'd91; b = 8'd225;  #10 
a = 8'd91; b = 8'd226;  #10 
a = 8'd91; b = 8'd227;  #10 
a = 8'd91; b = 8'd228;  #10 
a = 8'd91; b = 8'd229;  #10 
a = 8'd91; b = 8'd230;  #10 
a = 8'd91; b = 8'd231;  #10 
a = 8'd91; b = 8'd232;  #10 
a = 8'd91; b = 8'd233;  #10 
a = 8'd91; b = 8'd234;  #10 
a = 8'd91; b = 8'd235;  #10 
a = 8'd91; b = 8'd236;  #10 
a = 8'd91; b = 8'd237;  #10 
a = 8'd91; b = 8'd238;  #10 
a = 8'd91; b = 8'd239;  #10 
a = 8'd91; b = 8'd240;  #10 
a = 8'd91; b = 8'd241;  #10 
a = 8'd91; b = 8'd242;  #10 
a = 8'd91; b = 8'd243;  #10 
a = 8'd91; b = 8'd244;  #10 
a = 8'd91; b = 8'd245;  #10 
a = 8'd91; b = 8'd246;  #10 
a = 8'd91; b = 8'd247;  #10 
a = 8'd91; b = 8'd248;  #10 
a = 8'd91; b = 8'd249;  #10 
a = 8'd91; b = 8'd250;  #10 
a = 8'd91; b = 8'd251;  #10 
a = 8'd91; b = 8'd252;  #10 
a = 8'd91; b = 8'd253;  #10 
a = 8'd91; b = 8'd254;  #10 
a = 8'd91; b = 8'd255;  #10 
a = 8'd92; b = 8'd0;  #10 
a = 8'd92; b = 8'd1;  #10 
a = 8'd92; b = 8'd2;  #10 
a = 8'd92; b = 8'd3;  #10 
a = 8'd92; b = 8'd4;  #10 
a = 8'd92; b = 8'd5;  #10 
a = 8'd92; b = 8'd6;  #10 
a = 8'd92; b = 8'd7;  #10 
a = 8'd92; b = 8'd8;  #10 
a = 8'd92; b = 8'd9;  #10 
a = 8'd92; b = 8'd10;  #10 
a = 8'd92; b = 8'd11;  #10 
a = 8'd92; b = 8'd12;  #10 
a = 8'd92; b = 8'd13;  #10 
a = 8'd92; b = 8'd14;  #10 
a = 8'd92; b = 8'd15;  #10 
a = 8'd92; b = 8'd16;  #10 
a = 8'd92; b = 8'd17;  #10 
a = 8'd92; b = 8'd18;  #10 
a = 8'd92; b = 8'd19;  #10 
a = 8'd92; b = 8'd20;  #10 
a = 8'd92; b = 8'd21;  #10 
a = 8'd92; b = 8'd22;  #10 
a = 8'd92; b = 8'd23;  #10 
a = 8'd92; b = 8'd24;  #10 
a = 8'd92; b = 8'd25;  #10 
a = 8'd92; b = 8'd26;  #10 
a = 8'd92; b = 8'd27;  #10 
a = 8'd92; b = 8'd28;  #10 
a = 8'd92; b = 8'd29;  #10 
a = 8'd92; b = 8'd30;  #10 
a = 8'd92; b = 8'd31;  #10 
a = 8'd92; b = 8'd32;  #10 
a = 8'd92; b = 8'd33;  #10 
a = 8'd92; b = 8'd34;  #10 
a = 8'd92; b = 8'd35;  #10 
a = 8'd92; b = 8'd36;  #10 
a = 8'd92; b = 8'd37;  #10 
a = 8'd92; b = 8'd38;  #10 
a = 8'd92; b = 8'd39;  #10 
a = 8'd92; b = 8'd40;  #10 
a = 8'd92; b = 8'd41;  #10 
a = 8'd92; b = 8'd42;  #10 
a = 8'd92; b = 8'd43;  #10 
a = 8'd92; b = 8'd44;  #10 
a = 8'd92; b = 8'd45;  #10 
a = 8'd92; b = 8'd46;  #10 
a = 8'd92; b = 8'd47;  #10 
a = 8'd92; b = 8'd48;  #10 
a = 8'd92; b = 8'd49;  #10 
a = 8'd92; b = 8'd50;  #10 
a = 8'd92; b = 8'd51;  #10 
a = 8'd92; b = 8'd52;  #10 
a = 8'd92; b = 8'd53;  #10 
a = 8'd92; b = 8'd54;  #10 
a = 8'd92; b = 8'd55;  #10 
a = 8'd92; b = 8'd56;  #10 
a = 8'd92; b = 8'd57;  #10 
a = 8'd92; b = 8'd58;  #10 
a = 8'd92; b = 8'd59;  #10 
a = 8'd92; b = 8'd60;  #10 
a = 8'd92; b = 8'd61;  #10 
a = 8'd92; b = 8'd62;  #10 
a = 8'd92; b = 8'd63;  #10 
a = 8'd92; b = 8'd64;  #10 
a = 8'd92; b = 8'd65;  #10 
a = 8'd92; b = 8'd66;  #10 
a = 8'd92; b = 8'd67;  #10 
a = 8'd92; b = 8'd68;  #10 
a = 8'd92; b = 8'd69;  #10 
a = 8'd92; b = 8'd70;  #10 
a = 8'd92; b = 8'd71;  #10 
a = 8'd92; b = 8'd72;  #10 
a = 8'd92; b = 8'd73;  #10 
a = 8'd92; b = 8'd74;  #10 
a = 8'd92; b = 8'd75;  #10 
a = 8'd92; b = 8'd76;  #10 
a = 8'd92; b = 8'd77;  #10 
a = 8'd92; b = 8'd78;  #10 
a = 8'd92; b = 8'd79;  #10 
a = 8'd92; b = 8'd80;  #10 
a = 8'd92; b = 8'd81;  #10 
a = 8'd92; b = 8'd82;  #10 
a = 8'd92; b = 8'd83;  #10 
a = 8'd92; b = 8'd84;  #10 
a = 8'd92; b = 8'd85;  #10 
a = 8'd92; b = 8'd86;  #10 
a = 8'd92; b = 8'd87;  #10 
a = 8'd92; b = 8'd88;  #10 
a = 8'd92; b = 8'd89;  #10 
a = 8'd92; b = 8'd90;  #10 
a = 8'd92; b = 8'd91;  #10 
a = 8'd92; b = 8'd92;  #10 
a = 8'd92; b = 8'd93;  #10 
a = 8'd92; b = 8'd94;  #10 
a = 8'd92; b = 8'd95;  #10 
a = 8'd92; b = 8'd96;  #10 
a = 8'd92; b = 8'd97;  #10 
a = 8'd92; b = 8'd98;  #10 
a = 8'd92; b = 8'd99;  #10 
a = 8'd92; b = 8'd100;  #10 
a = 8'd92; b = 8'd101;  #10 
a = 8'd92; b = 8'd102;  #10 
a = 8'd92; b = 8'd103;  #10 
a = 8'd92; b = 8'd104;  #10 
a = 8'd92; b = 8'd105;  #10 
a = 8'd92; b = 8'd106;  #10 
a = 8'd92; b = 8'd107;  #10 
a = 8'd92; b = 8'd108;  #10 
a = 8'd92; b = 8'd109;  #10 
a = 8'd92; b = 8'd110;  #10 
a = 8'd92; b = 8'd111;  #10 
a = 8'd92; b = 8'd112;  #10 
a = 8'd92; b = 8'd113;  #10 
a = 8'd92; b = 8'd114;  #10 
a = 8'd92; b = 8'd115;  #10 
a = 8'd92; b = 8'd116;  #10 
a = 8'd92; b = 8'd117;  #10 
a = 8'd92; b = 8'd118;  #10 
a = 8'd92; b = 8'd119;  #10 
a = 8'd92; b = 8'd120;  #10 
a = 8'd92; b = 8'd121;  #10 
a = 8'd92; b = 8'd122;  #10 
a = 8'd92; b = 8'd123;  #10 
a = 8'd92; b = 8'd124;  #10 
a = 8'd92; b = 8'd125;  #10 
a = 8'd92; b = 8'd126;  #10 
a = 8'd92; b = 8'd127;  #10 
a = 8'd92; b = 8'd128;  #10 
a = 8'd92; b = 8'd129;  #10 
a = 8'd92; b = 8'd130;  #10 
a = 8'd92; b = 8'd131;  #10 
a = 8'd92; b = 8'd132;  #10 
a = 8'd92; b = 8'd133;  #10 
a = 8'd92; b = 8'd134;  #10 
a = 8'd92; b = 8'd135;  #10 
a = 8'd92; b = 8'd136;  #10 
a = 8'd92; b = 8'd137;  #10 
a = 8'd92; b = 8'd138;  #10 
a = 8'd92; b = 8'd139;  #10 
a = 8'd92; b = 8'd140;  #10 
a = 8'd92; b = 8'd141;  #10 
a = 8'd92; b = 8'd142;  #10 
a = 8'd92; b = 8'd143;  #10 
a = 8'd92; b = 8'd144;  #10 
a = 8'd92; b = 8'd145;  #10 
a = 8'd92; b = 8'd146;  #10 
a = 8'd92; b = 8'd147;  #10 
a = 8'd92; b = 8'd148;  #10 
a = 8'd92; b = 8'd149;  #10 
a = 8'd92; b = 8'd150;  #10 
a = 8'd92; b = 8'd151;  #10 
a = 8'd92; b = 8'd152;  #10 
a = 8'd92; b = 8'd153;  #10 
a = 8'd92; b = 8'd154;  #10 
a = 8'd92; b = 8'd155;  #10 
a = 8'd92; b = 8'd156;  #10 
a = 8'd92; b = 8'd157;  #10 
a = 8'd92; b = 8'd158;  #10 
a = 8'd92; b = 8'd159;  #10 
a = 8'd92; b = 8'd160;  #10 
a = 8'd92; b = 8'd161;  #10 
a = 8'd92; b = 8'd162;  #10 
a = 8'd92; b = 8'd163;  #10 
a = 8'd92; b = 8'd164;  #10 
a = 8'd92; b = 8'd165;  #10 
a = 8'd92; b = 8'd166;  #10 
a = 8'd92; b = 8'd167;  #10 
a = 8'd92; b = 8'd168;  #10 
a = 8'd92; b = 8'd169;  #10 
a = 8'd92; b = 8'd170;  #10 
a = 8'd92; b = 8'd171;  #10 
a = 8'd92; b = 8'd172;  #10 
a = 8'd92; b = 8'd173;  #10 
a = 8'd92; b = 8'd174;  #10 
a = 8'd92; b = 8'd175;  #10 
a = 8'd92; b = 8'd176;  #10 
a = 8'd92; b = 8'd177;  #10 
a = 8'd92; b = 8'd178;  #10 
a = 8'd92; b = 8'd179;  #10 
a = 8'd92; b = 8'd180;  #10 
a = 8'd92; b = 8'd181;  #10 
a = 8'd92; b = 8'd182;  #10 
a = 8'd92; b = 8'd183;  #10 
a = 8'd92; b = 8'd184;  #10 
a = 8'd92; b = 8'd185;  #10 
a = 8'd92; b = 8'd186;  #10 
a = 8'd92; b = 8'd187;  #10 
a = 8'd92; b = 8'd188;  #10 
a = 8'd92; b = 8'd189;  #10 
a = 8'd92; b = 8'd190;  #10 
a = 8'd92; b = 8'd191;  #10 
a = 8'd92; b = 8'd192;  #10 
a = 8'd92; b = 8'd193;  #10 
a = 8'd92; b = 8'd194;  #10 
a = 8'd92; b = 8'd195;  #10 
a = 8'd92; b = 8'd196;  #10 
a = 8'd92; b = 8'd197;  #10 
a = 8'd92; b = 8'd198;  #10 
a = 8'd92; b = 8'd199;  #10 
a = 8'd92; b = 8'd200;  #10 
a = 8'd92; b = 8'd201;  #10 
a = 8'd92; b = 8'd202;  #10 
a = 8'd92; b = 8'd203;  #10 
a = 8'd92; b = 8'd204;  #10 
a = 8'd92; b = 8'd205;  #10 
a = 8'd92; b = 8'd206;  #10 
a = 8'd92; b = 8'd207;  #10 
a = 8'd92; b = 8'd208;  #10 
a = 8'd92; b = 8'd209;  #10 
a = 8'd92; b = 8'd210;  #10 
a = 8'd92; b = 8'd211;  #10 
a = 8'd92; b = 8'd212;  #10 
a = 8'd92; b = 8'd213;  #10 
a = 8'd92; b = 8'd214;  #10 
a = 8'd92; b = 8'd215;  #10 
a = 8'd92; b = 8'd216;  #10 
a = 8'd92; b = 8'd217;  #10 
a = 8'd92; b = 8'd218;  #10 
a = 8'd92; b = 8'd219;  #10 
a = 8'd92; b = 8'd220;  #10 
a = 8'd92; b = 8'd221;  #10 
a = 8'd92; b = 8'd222;  #10 
a = 8'd92; b = 8'd223;  #10 
a = 8'd92; b = 8'd224;  #10 
a = 8'd92; b = 8'd225;  #10 
a = 8'd92; b = 8'd226;  #10 
a = 8'd92; b = 8'd227;  #10 
a = 8'd92; b = 8'd228;  #10 
a = 8'd92; b = 8'd229;  #10 
a = 8'd92; b = 8'd230;  #10 
a = 8'd92; b = 8'd231;  #10 
a = 8'd92; b = 8'd232;  #10 
a = 8'd92; b = 8'd233;  #10 
a = 8'd92; b = 8'd234;  #10 
a = 8'd92; b = 8'd235;  #10 
a = 8'd92; b = 8'd236;  #10 
a = 8'd92; b = 8'd237;  #10 
a = 8'd92; b = 8'd238;  #10 
a = 8'd92; b = 8'd239;  #10 
a = 8'd92; b = 8'd240;  #10 
a = 8'd92; b = 8'd241;  #10 
a = 8'd92; b = 8'd242;  #10 
a = 8'd92; b = 8'd243;  #10 
a = 8'd92; b = 8'd244;  #10 
a = 8'd92; b = 8'd245;  #10 
a = 8'd92; b = 8'd246;  #10 
a = 8'd92; b = 8'd247;  #10 
a = 8'd92; b = 8'd248;  #10 
a = 8'd92; b = 8'd249;  #10 
a = 8'd92; b = 8'd250;  #10 
a = 8'd92; b = 8'd251;  #10 
a = 8'd92; b = 8'd252;  #10 
a = 8'd92; b = 8'd253;  #10 
a = 8'd92; b = 8'd254;  #10 
a = 8'd92; b = 8'd255;  #10 
a = 8'd93; b = 8'd0;  #10 
a = 8'd93; b = 8'd1;  #10 
a = 8'd93; b = 8'd2;  #10 
a = 8'd93; b = 8'd3;  #10 
a = 8'd93; b = 8'd4;  #10 
a = 8'd93; b = 8'd5;  #10 
a = 8'd93; b = 8'd6;  #10 
a = 8'd93; b = 8'd7;  #10 
a = 8'd93; b = 8'd8;  #10 
a = 8'd93; b = 8'd9;  #10 
a = 8'd93; b = 8'd10;  #10 
a = 8'd93; b = 8'd11;  #10 
a = 8'd93; b = 8'd12;  #10 
a = 8'd93; b = 8'd13;  #10 
a = 8'd93; b = 8'd14;  #10 
a = 8'd93; b = 8'd15;  #10 
a = 8'd93; b = 8'd16;  #10 
a = 8'd93; b = 8'd17;  #10 
a = 8'd93; b = 8'd18;  #10 
a = 8'd93; b = 8'd19;  #10 
a = 8'd93; b = 8'd20;  #10 
a = 8'd93; b = 8'd21;  #10 
a = 8'd93; b = 8'd22;  #10 
a = 8'd93; b = 8'd23;  #10 
a = 8'd93; b = 8'd24;  #10 
a = 8'd93; b = 8'd25;  #10 
a = 8'd93; b = 8'd26;  #10 
a = 8'd93; b = 8'd27;  #10 
a = 8'd93; b = 8'd28;  #10 
a = 8'd93; b = 8'd29;  #10 
a = 8'd93; b = 8'd30;  #10 
a = 8'd93; b = 8'd31;  #10 
a = 8'd93; b = 8'd32;  #10 
a = 8'd93; b = 8'd33;  #10 
a = 8'd93; b = 8'd34;  #10 
a = 8'd93; b = 8'd35;  #10 
a = 8'd93; b = 8'd36;  #10 
a = 8'd93; b = 8'd37;  #10 
a = 8'd93; b = 8'd38;  #10 
a = 8'd93; b = 8'd39;  #10 
a = 8'd93; b = 8'd40;  #10 
a = 8'd93; b = 8'd41;  #10 
a = 8'd93; b = 8'd42;  #10 
a = 8'd93; b = 8'd43;  #10 
a = 8'd93; b = 8'd44;  #10 
a = 8'd93; b = 8'd45;  #10 
a = 8'd93; b = 8'd46;  #10 
a = 8'd93; b = 8'd47;  #10 
a = 8'd93; b = 8'd48;  #10 
a = 8'd93; b = 8'd49;  #10 
a = 8'd93; b = 8'd50;  #10 
a = 8'd93; b = 8'd51;  #10 
a = 8'd93; b = 8'd52;  #10 
a = 8'd93; b = 8'd53;  #10 
a = 8'd93; b = 8'd54;  #10 
a = 8'd93; b = 8'd55;  #10 
a = 8'd93; b = 8'd56;  #10 
a = 8'd93; b = 8'd57;  #10 
a = 8'd93; b = 8'd58;  #10 
a = 8'd93; b = 8'd59;  #10 
a = 8'd93; b = 8'd60;  #10 
a = 8'd93; b = 8'd61;  #10 
a = 8'd93; b = 8'd62;  #10 
a = 8'd93; b = 8'd63;  #10 
a = 8'd93; b = 8'd64;  #10 
a = 8'd93; b = 8'd65;  #10 
a = 8'd93; b = 8'd66;  #10 
a = 8'd93; b = 8'd67;  #10 
a = 8'd93; b = 8'd68;  #10 
a = 8'd93; b = 8'd69;  #10 
a = 8'd93; b = 8'd70;  #10 
a = 8'd93; b = 8'd71;  #10 
a = 8'd93; b = 8'd72;  #10 
a = 8'd93; b = 8'd73;  #10 
a = 8'd93; b = 8'd74;  #10 
a = 8'd93; b = 8'd75;  #10 
a = 8'd93; b = 8'd76;  #10 
a = 8'd93; b = 8'd77;  #10 
a = 8'd93; b = 8'd78;  #10 
a = 8'd93; b = 8'd79;  #10 
a = 8'd93; b = 8'd80;  #10 
a = 8'd93; b = 8'd81;  #10 
a = 8'd93; b = 8'd82;  #10 
a = 8'd93; b = 8'd83;  #10 
a = 8'd93; b = 8'd84;  #10 
a = 8'd93; b = 8'd85;  #10 
a = 8'd93; b = 8'd86;  #10 
a = 8'd93; b = 8'd87;  #10 
a = 8'd93; b = 8'd88;  #10 
a = 8'd93; b = 8'd89;  #10 
a = 8'd93; b = 8'd90;  #10 
a = 8'd93; b = 8'd91;  #10 
a = 8'd93; b = 8'd92;  #10 
a = 8'd93; b = 8'd93;  #10 
a = 8'd93; b = 8'd94;  #10 
a = 8'd93; b = 8'd95;  #10 
a = 8'd93; b = 8'd96;  #10 
a = 8'd93; b = 8'd97;  #10 
a = 8'd93; b = 8'd98;  #10 
a = 8'd93; b = 8'd99;  #10 
a = 8'd93; b = 8'd100;  #10 
a = 8'd93; b = 8'd101;  #10 
a = 8'd93; b = 8'd102;  #10 
a = 8'd93; b = 8'd103;  #10 
a = 8'd93; b = 8'd104;  #10 
a = 8'd93; b = 8'd105;  #10 
a = 8'd93; b = 8'd106;  #10 
a = 8'd93; b = 8'd107;  #10 
a = 8'd93; b = 8'd108;  #10 
a = 8'd93; b = 8'd109;  #10 
a = 8'd93; b = 8'd110;  #10 
a = 8'd93; b = 8'd111;  #10 
a = 8'd93; b = 8'd112;  #10 
a = 8'd93; b = 8'd113;  #10 
a = 8'd93; b = 8'd114;  #10 
a = 8'd93; b = 8'd115;  #10 
a = 8'd93; b = 8'd116;  #10 
a = 8'd93; b = 8'd117;  #10 
a = 8'd93; b = 8'd118;  #10 
a = 8'd93; b = 8'd119;  #10 
a = 8'd93; b = 8'd120;  #10 
a = 8'd93; b = 8'd121;  #10 
a = 8'd93; b = 8'd122;  #10 
a = 8'd93; b = 8'd123;  #10 
a = 8'd93; b = 8'd124;  #10 
a = 8'd93; b = 8'd125;  #10 
a = 8'd93; b = 8'd126;  #10 
a = 8'd93; b = 8'd127;  #10 
a = 8'd93; b = 8'd128;  #10 
a = 8'd93; b = 8'd129;  #10 
a = 8'd93; b = 8'd130;  #10 
a = 8'd93; b = 8'd131;  #10 
a = 8'd93; b = 8'd132;  #10 
a = 8'd93; b = 8'd133;  #10 
a = 8'd93; b = 8'd134;  #10 
a = 8'd93; b = 8'd135;  #10 
a = 8'd93; b = 8'd136;  #10 
a = 8'd93; b = 8'd137;  #10 
a = 8'd93; b = 8'd138;  #10 
a = 8'd93; b = 8'd139;  #10 
a = 8'd93; b = 8'd140;  #10 
a = 8'd93; b = 8'd141;  #10 
a = 8'd93; b = 8'd142;  #10 
a = 8'd93; b = 8'd143;  #10 
a = 8'd93; b = 8'd144;  #10 
a = 8'd93; b = 8'd145;  #10 
a = 8'd93; b = 8'd146;  #10 
a = 8'd93; b = 8'd147;  #10 
a = 8'd93; b = 8'd148;  #10 
a = 8'd93; b = 8'd149;  #10 
a = 8'd93; b = 8'd150;  #10 
a = 8'd93; b = 8'd151;  #10 
a = 8'd93; b = 8'd152;  #10 
a = 8'd93; b = 8'd153;  #10 
a = 8'd93; b = 8'd154;  #10 
a = 8'd93; b = 8'd155;  #10 
a = 8'd93; b = 8'd156;  #10 
a = 8'd93; b = 8'd157;  #10 
a = 8'd93; b = 8'd158;  #10 
a = 8'd93; b = 8'd159;  #10 
a = 8'd93; b = 8'd160;  #10 
a = 8'd93; b = 8'd161;  #10 
a = 8'd93; b = 8'd162;  #10 
a = 8'd93; b = 8'd163;  #10 
a = 8'd93; b = 8'd164;  #10 
a = 8'd93; b = 8'd165;  #10 
a = 8'd93; b = 8'd166;  #10 
a = 8'd93; b = 8'd167;  #10 
a = 8'd93; b = 8'd168;  #10 
a = 8'd93; b = 8'd169;  #10 
a = 8'd93; b = 8'd170;  #10 
a = 8'd93; b = 8'd171;  #10 
a = 8'd93; b = 8'd172;  #10 
a = 8'd93; b = 8'd173;  #10 
a = 8'd93; b = 8'd174;  #10 
a = 8'd93; b = 8'd175;  #10 
a = 8'd93; b = 8'd176;  #10 
a = 8'd93; b = 8'd177;  #10 
a = 8'd93; b = 8'd178;  #10 
a = 8'd93; b = 8'd179;  #10 
a = 8'd93; b = 8'd180;  #10 
a = 8'd93; b = 8'd181;  #10 
a = 8'd93; b = 8'd182;  #10 
a = 8'd93; b = 8'd183;  #10 
a = 8'd93; b = 8'd184;  #10 
a = 8'd93; b = 8'd185;  #10 
a = 8'd93; b = 8'd186;  #10 
a = 8'd93; b = 8'd187;  #10 
a = 8'd93; b = 8'd188;  #10 
a = 8'd93; b = 8'd189;  #10 
a = 8'd93; b = 8'd190;  #10 
a = 8'd93; b = 8'd191;  #10 
a = 8'd93; b = 8'd192;  #10 
a = 8'd93; b = 8'd193;  #10 
a = 8'd93; b = 8'd194;  #10 
a = 8'd93; b = 8'd195;  #10 
a = 8'd93; b = 8'd196;  #10 
a = 8'd93; b = 8'd197;  #10 
a = 8'd93; b = 8'd198;  #10 
a = 8'd93; b = 8'd199;  #10 
a = 8'd93; b = 8'd200;  #10 
a = 8'd93; b = 8'd201;  #10 
a = 8'd93; b = 8'd202;  #10 
a = 8'd93; b = 8'd203;  #10 
a = 8'd93; b = 8'd204;  #10 
a = 8'd93; b = 8'd205;  #10 
a = 8'd93; b = 8'd206;  #10 
a = 8'd93; b = 8'd207;  #10 
a = 8'd93; b = 8'd208;  #10 
a = 8'd93; b = 8'd209;  #10 
a = 8'd93; b = 8'd210;  #10 
a = 8'd93; b = 8'd211;  #10 
a = 8'd93; b = 8'd212;  #10 
a = 8'd93; b = 8'd213;  #10 
a = 8'd93; b = 8'd214;  #10 
a = 8'd93; b = 8'd215;  #10 
a = 8'd93; b = 8'd216;  #10 
a = 8'd93; b = 8'd217;  #10 
a = 8'd93; b = 8'd218;  #10 
a = 8'd93; b = 8'd219;  #10 
a = 8'd93; b = 8'd220;  #10 
a = 8'd93; b = 8'd221;  #10 
a = 8'd93; b = 8'd222;  #10 
a = 8'd93; b = 8'd223;  #10 
a = 8'd93; b = 8'd224;  #10 
a = 8'd93; b = 8'd225;  #10 
a = 8'd93; b = 8'd226;  #10 
a = 8'd93; b = 8'd227;  #10 
a = 8'd93; b = 8'd228;  #10 
a = 8'd93; b = 8'd229;  #10 
a = 8'd93; b = 8'd230;  #10 
a = 8'd93; b = 8'd231;  #10 
a = 8'd93; b = 8'd232;  #10 
a = 8'd93; b = 8'd233;  #10 
a = 8'd93; b = 8'd234;  #10 
a = 8'd93; b = 8'd235;  #10 
a = 8'd93; b = 8'd236;  #10 
a = 8'd93; b = 8'd237;  #10 
a = 8'd93; b = 8'd238;  #10 
a = 8'd93; b = 8'd239;  #10 
a = 8'd93; b = 8'd240;  #10 
a = 8'd93; b = 8'd241;  #10 
a = 8'd93; b = 8'd242;  #10 
a = 8'd93; b = 8'd243;  #10 
a = 8'd93; b = 8'd244;  #10 
a = 8'd93; b = 8'd245;  #10 
a = 8'd93; b = 8'd246;  #10 
a = 8'd93; b = 8'd247;  #10 
a = 8'd93; b = 8'd248;  #10 
a = 8'd93; b = 8'd249;  #10 
a = 8'd93; b = 8'd250;  #10 
a = 8'd93; b = 8'd251;  #10 
a = 8'd93; b = 8'd252;  #10 
a = 8'd93; b = 8'd253;  #10 
a = 8'd93; b = 8'd254;  #10 
a = 8'd93; b = 8'd255;  #10 
a = 8'd94; b = 8'd0;  #10 
a = 8'd94; b = 8'd1;  #10 
a = 8'd94; b = 8'd2;  #10 
a = 8'd94; b = 8'd3;  #10 
a = 8'd94; b = 8'd4;  #10 
a = 8'd94; b = 8'd5;  #10 
a = 8'd94; b = 8'd6;  #10 
a = 8'd94; b = 8'd7;  #10 
a = 8'd94; b = 8'd8;  #10 
a = 8'd94; b = 8'd9;  #10 
a = 8'd94; b = 8'd10;  #10 
a = 8'd94; b = 8'd11;  #10 
a = 8'd94; b = 8'd12;  #10 
a = 8'd94; b = 8'd13;  #10 
a = 8'd94; b = 8'd14;  #10 
a = 8'd94; b = 8'd15;  #10 
a = 8'd94; b = 8'd16;  #10 
a = 8'd94; b = 8'd17;  #10 
a = 8'd94; b = 8'd18;  #10 
a = 8'd94; b = 8'd19;  #10 
a = 8'd94; b = 8'd20;  #10 
a = 8'd94; b = 8'd21;  #10 
a = 8'd94; b = 8'd22;  #10 
a = 8'd94; b = 8'd23;  #10 
a = 8'd94; b = 8'd24;  #10 
a = 8'd94; b = 8'd25;  #10 
a = 8'd94; b = 8'd26;  #10 
a = 8'd94; b = 8'd27;  #10 
a = 8'd94; b = 8'd28;  #10 
a = 8'd94; b = 8'd29;  #10 
a = 8'd94; b = 8'd30;  #10 
a = 8'd94; b = 8'd31;  #10 
a = 8'd94; b = 8'd32;  #10 
a = 8'd94; b = 8'd33;  #10 
a = 8'd94; b = 8'd34;  #10 
a = 8'd94; b = 8'd35;  #10 
a = 8'd94; b = 8'd36;  #10 
a = 8'd94; b = 8'd37;  #10 
a = 8'd94; b = 8'd38;  #10 
a = 8'd94; b = 8'd39;  #10 
a = 8'd94; b = 8'd40;  #10 
a = 8'd94; b = 8'd41;  #10 
a = 8'd94; b = 8'd42;  #10 
a = 8'd94; b = 8'd43;  #10 
a = 8'd94; b = 8'd44;  #10 
a = 8'd94; b = 8'd45;  #10 
a = 8'd94; b = 8'd46;  #10 
a = 8'd94; b = 8'd47;  #10 
a = 8'd94; b = 8'd48;  #10 
a = 8'd94; b = 8'd49;  #10 
a = 8'd94; b = 8'd50;  #10 
a = 8'd94; b = 8'd51;  #10 
a = 8'd94; b = 8'd52;  #10 
a = 8'd94; b = 8'd53;  #10 
a = 8'd94; b = 8'd54;  #10 
a = 8'd94; b = 8'd55;  #10 
a = 8'd94; b = 8'd56;  #10 
a = 8'd94; b = 8'd57;  #10 
a = 8'd94; b = 8'd58;  #10 
a = 8'd94; b = 8'd59;  #10 
a = 8'd94; b = 8'd60;  #10 
a = 8'd94; b = 8'd61;  #10 
a = 8'd94; b = 8'd62;  #10 
a = 8'd94; b = 8'd63;  #10 
a = 8'd94; b = 8'd64;  #10 
a = 8'd94; b = 8'd65;  #10 
a = 8'd94; b = 8'd66;  #10 
a = 8'd94; b = 8'd67;  #10 
a = 8'd94; b = 8'd68;  #10 
a = 8'd94; b = 8'd69;  #10 
a = 8'd94; b = 8'd70;  #10 
a = 8'd94; b = 8'd71;  #10 
a = 8'd94; b = 8'd72;  #10 
a = 8'd94; b = 8'd73;  #10 
a = 8'd94; b = 8'd74;  #10 
a = 8'd94; b = 8'd75;  #10 
a = 8'd94; b = 8'd76;  #10 
a = 8'd94; b = 8'd77;  #10 
a = 8'd94; b = 8'd78;  #10 
a = 8'd94; b = 8'd79;  #10 
a = 8'd94; b = 8'd80;  #10 
a = 8'd94; b = 8'd81;  #10 
a = 8'd94; b = 8'd82;  #10 
a = 8'd94; b = 8'd83;  #10 
a = 8'd94; b = 8'd84;  #10 
a = 8'd94; b = 8'd85;  #10 
a = 8'd94; b = 8'd86;  #10 
a = 8'd94; b = 8'd87;  #10 
a = 8'd94; b = 8'd88;  #10 
a = 8'd94; b = 8'd89;  #10 
a = 8'd94; b = 8'd90;  #10 
a = 8'd94; b = 8'd91;  #10 
a = 8'd94; b = 8'd92;  #10 
a = 8'd94; b = 8'd93;  #10 
a = 8'd94; b = 8'd94;  #10 
a = 8'd94; b = 8'd95;  #10 
a = 8'd94; b = 8'd96;  #10 
a = 8'd94; b = 8'd97;  #10 
a = 8'd94; b = 8'd98;  #10 
a = 8'd94; b = 8'd99;  #10 
a = 8'd94; b = 8'd100;  #10 
a = 8'd94; b = 8'd101;  #10 
a = 8'd94; b = 8'd102;  #10 
a = 8'd94; b = 8'd103;  #10 
a = 8'd94; b = 8'd104;  #10 
a = 8'd94; b = 8'd105;  #10 
a = 8'd94; b = 8'd106;  #10 
a = 8'd94; b = 8'd107;  #10 
a = 8'd94; b = 8'd108;  #10 
a = 8'd94; b = 8'd109;  #10 
a = 8'd94; b = 8'd110;  #10 
a = 8'd94; b = 8'd111;  #10 
a = 8'd94; b = 8'd112;  #10 
a = 8'd94; b = 8'd113;  #10 
a = 8'd94; b = 8'd114;  #10 
a = 8'd94; b = 8'd115;  #10 
a = 8'd94; b = 8'd116;  #10 
a = 8'd94; b = 8'd117;  #10 
a = 8'd94; b = 8'd118;  #10 
a = 8'd94; b = 8'd119;  #10 
a = 8'd94; b = 8'd120;  #10 
a = 8'd94; b = 8'd121;  #10 
a = 8'd94; b = 8'd122;  #10 
a = 8'd94; b = 8'd123;  #10 
a = 8'd94; b = 8'd124;  #10 
a = 8'd94; b = 8'd125;  #10 
a = 8'd94; b = 8'd126;  #10 
a = 8'd94; b = 8'd127;  #10 
a = 8'd94; b = 8'd128;  #10 
a = 8'd94; b = 8'd129;  #10 
a = 8'd94; b = 8'd130;  #10 
a = 8'd94; b = 8'd131;  #10 
a = 8'd94; b = 8'd132;  #10 
a = 8'd94; b = 8'd133;  #10 
a = 8'd94; b = 8'd134;  #10 
a = 8'd94; b = 8'd135;  #10 
a = 8'd94; b = 8'd136;  #10 
a = 8'd94; b = 8'd137;  #10 
a = 8'd94; b = 8'd138;  #10 
a = 8'd94; b = 8'd139;  #10 
a = 8'd94; b = 8'd140;  #10 
a = 8'd94; b = 8'd141;  #10 
a = 8'd94; b = 8'd142;  #10 
a = 8'd94; b = 8'd143;  #10 
a = 8'd94; b = 8'd144;  #10 
a = 8'd94; b = 8'd145;  #10 
a = 8'd94; b = 8'd146;  #10 
a = 8'd94; b = 8'd147;  #10 
a = 8'd94; b = 8'd148;  #10 
a = 8'd94; b = 8'd149;  #10 
a = 8'd94; b = 8'd150;  #10 
a = 8'd94; b = 8'd151;  #10 
a = 8'd94; b = 8'd152;  #10 
a = 8'd94; b = 8'd153;  #10 
a = 8'd94; b = 8'd154;  #10 
a = 8'd94; b = 8'd155;  #10 
a = 8'd94; b = 8'd156;  #10 
a = 8'd94; b = 8'd157;  #10 
a = 8'd94; b = 8'd158;  #10 
a = 8'd94; b = 8'd159;  #10 
a = 8'd94; b = 8'd160;  #10 
a = 8'd94; b = 8'd161;  #10 
a = 8'd94; b = 8'd162;  #10 
a = 8'd94; b = 8'd163;  #10 
a = 8'd94; b = 8'd164;  #10 
a = 8'd94; b = 8'd165;  #10 
a = 8'd94; b = 8'd166;  #10 
a = 8'd94; b = 8'd167;  #10 
a = 8'd94; b = 8'd168;  #10 
a = 8'd94; b = 8'd169;  #10 
a = 8'd94; b = 8'd170;  #10 
a = 8'd94; b = 8'd171;  #10 
a = 8'd94; b = 8'd172;  #10 
a = 8'd94; b = 8'd173;  #10 
a = 8'd94; b = 8'd174;  #10 
a = 8'd94; b = 8'd175;  #10 
a = 8'd94; b = 8'd176;  #10 
a = 8'd94; b = 8'd177;  #10 
a = 8'd94; b = 8'd178;  #10 
a = 8'd94; b = 8'd179;  #10 
a = 8'd94; b = 8'd180;  #10 
a = 8'd94; b = 8'd181;  #10 
a = 8'd94; b = 8'd182;  #10 
a = 8'd94; b = 8'd183;  #10 
a = 8'd94; b = 8'd184;  #10 
a = 8'd94; b = 8'd185;  #10 
a = 8'd94; b = 8'd186;  #10 
a = 8'd94; b = 8'd187;  #10 
a = 8'd94; b = 8'd188;  #10 
a = 8'd94; b = 8'd189;  #10 
a = 8'd94; b = 8'd190;  #10 
a = 8'd94; b = 8'd191;  #10 
a = 8'd94; b = 8'd192;  #10 
a = 8'd94; b = 8'd193;  #10 
a = 8'd94; b = 8'd194;  #10 
a = 8'd94; b = 8'd195;  #10 
a = 8'd94; b = 8'd196;  #10 
a = 8'd94; b = 8'd197;  #10 
a = 8'd94; b = 8'd198;  #10 
a = 8'd94; b = 8'd199;  #10 
a = 8'd94; b = 8'd200;  #10 
a = 8'd94; b = 8'd201;  #10 
a = 8'd94; b = 8'd202;  #10 
a = 8'd94; b = 8'd203;  #10 
a = 8'd94; b = 8'd204;  #10 
a = 8'd94; b = 8'd205;  #10 
a = 8'd94; b = 8'd206;  #10 
a = 8'd94; b = 8'd207;  #10 
a = 8'd94; b = 8'd208;  #10 
a = 8'd94; b = 8'd209;  #10 
a = 8'd94; b = 8'd210;  #10 
a = 8'd94; b = 8'd211;  #10 
a = 8'd94; b = 8'd212;  #10 
a = 8'd94; b = 8'd213;  #10 
a = 8'd94; b = 8'd214;  #10 
a = 8'd94; b = 8'd215;  #10 
a = 8'd94; b = 8'd216;  #10 
a = 8'd94; b = 8'd217;  #10 
a = 8'd94; b = 8'd218;  #10 
a = 8'd94; b = 8'd219;  #10 
a = 8'd94; b = 8'd220;  #10 
a = 8'd94; b = 8'd221;  #10 
a = 8'd94; b = 8'd222;  #10 
a = 8'd94; b = 8'd223;  #10 
a = 8'd94; b = 8'd224;  #10 
a = 8'd94; b = 8'd225;  #10 
a = 8'd94; b = 8'd226;  #10 
a = 8'd94; b = 8'd227;  #10 
a = 8'd94; b = 8'd228;  #10 
a = 8'd94; b = 8'd229;  #10 
a = 8'd94; b = 8'd230;  #10 
a = 8'd94; b = 8'd231;  #10 
a = 8'd94; b = 8'd232;  #10 
a = 8'd94; b = 8'd233;  #10 
a = 8'd94; b = 8'd234;  #10 
a = 8'd94; b = 8'd235;  #10 
a = 8'd94; b = 8'd236;  #10 
a = 8'd94; b = 8'd237;  #10 
a = 8'd94; b = 8'd238;  #10 
a = 8'd94; b = 8'd239;  #10 
a = 8'd94; b = 8'd240;  #10 
a = 8'd94; b = 8'd241;  #10 
a = 8'd94; b = 8'd242;  #10 
a = 8'd94; b = 8'd243;  #10 
a = 8'd94; b = 8'd244;  #10 
a = 8'd94; b = 8'd245;  #10 
a = 8'd94; b = 8'd246;  #10 
a = 8'd94; b = 8'd247;  #10 
a = 8'd94; b = 8'd248;  #10 
a = 8'd94; b = 8'd249;  #10 
a = 8'd94; b = 8'd250;  #10 
a = 8'd94; b = 8'd251;  #10 
a = 8'd94; b = 8'd252;  #10 
a = 8'd94; b = 8'd253;  #10 
a = 8'd94; b = 8'd254;  #10 
a = 8'd94; b = 8'd255;  #10 
a = 8'd95; b = 8'd0;  #10 
a = 8'd95; b = 8'd1;  #10 
a = 8'd95; b = 8'd2;  #10 
a = 8'd95; b = 8'd3;  #10 
a = 8'd95; b = 8'd4;  #10 
a = 8'd95; b = 8'd5;  #10 
a = 8'd95; b = 8'd6;  #10 
a = 8'd95; b = 8'd7;  #10 
a = 8'd95; b = 8'd8;  #10 
a = 8'd95; b = 8'd9;  #10 
a = 8'd95; b = 8'd10;  #10 
a = 8'd95; b = 8'd11;  #10 
a = 8'd95; b = 8'd12;  #10 
a = 8'd95; b = 8'd13;  #10 
a = 8'd95; b = 8'd14;  #10 
a = 8'd95; b = 8'd15;  #10 
a = 8'd95; b = 8'd16;  #10 
a = 8'd95; b = 8'd17;  #10 
a = 8'd95; b = 8'd18;  #10 
a = 8'd95; b = 8'd19;  #10 
a = 8'd95; b = 8'd20;  #10 
a = 8'd95; b = 8'd21;  #10 
a = 8'd95; b = 8'd22;  #10 
a = 8'd95; b = 8'd23;  #10 
a = 8'd95; b = 8'd24;  #10 
a = 8'd95; b = 8'd25;  #10 
a = 8'd95; b = 8'd26;  #10 
a = 8'd95; b = 8'd27;  #10 
a = 8'd95; b = 8'd28;  #10 
a = 8'd95; b = 8'd29;  #10 
a = 8'd95; b = 8'd30;  #10 
a = 8'd95; b = 8'd31;  #10 
a = 8'd95; b = 8'd32;  #10 
a = 8'd95; b = 8'd33;  #10 
a = 8'd95; b = 8'd34;  #10 
a = 8'd95; b = 8'd35;  #10 
a = 8'd95; b = 8'd36;  #10 
a = 8'd95; b = 8'd37;  #10 
a = 8'd95; b = 8'd38;  #10 
a = 8'd95; b = 8'd39;  #10 
a = 8'd95; b = 8'd40;  #10 
a = 8'd95; b = 8'd41;  #10 
a = 8'd95; b = 8'd42;  #10 
a = 8'd95; b = 8'd43;  #10 
a = 8'd95; b = 8'd44;  #10 
a = 8'd95; b = 8'd45;  #10 
a = 8'd95; b = 8'd46;  #10 
a = 8'd95; b = 8'd47;  #10 
a = 8'd95; b = 8'd48;  #10 
a = 8'd95; b = 8'd49;  #10 
a = 8'd95; b = 8'd50;  #10 
a = 8'd95; b = 8'd51;  #10 
a = 8'd95; b = 8'd52;  #10 
a = 8'd95; b = 8'd53;  #10 
a = 8'd95; b = 8'd54;  #10 
a = 8'd95; b = 8'd55;  #10 
a = 8'd95; b = 8'd56;  #10 
a = 8'd95; b = 8'd57;  #10 
a = 8'd95; b = 8'd58;  #10 
a = 8'd95; b = 8'd59;  #10 
a = 8'd95; b = 8'd60;  #10 
a = 8'd95; b = 8'd61;  #10 
a = 8'd95; b = 8'd62;  #10 
a = 8'd95; b = 8'd63;  #10 
a = 8'd95; b = 8'd64;  #10 
a = 8'd95; b = 8'd65;  #10 
a = 8'd95; b = 8'd66;  #10 
a = 8'd95; b = 8'd67;  #10 
a = 8'd95; b = 8'd68;  #10 
a = 8'd95; b = 8'd69;  #10 
a = 8'd95; b = 8'd70;  #10 
a = 8'd95; b = 8'd71;  #10 
a = 8'd95; b = 8'd72;  #10 
a = 8'd95; b = 8'd73;  #10 
a = 8'd95; b = 8'd74;  #10 
a = 8'd95; b = 8'd75;  #10 
a = 8'd95; b = 8'd76;  #10 
a = 8'd95; b = 8'd77;  #10 
a = 8'd95; b = 8'd78;  #10 
a = 8'd95; b = 8'd79;  #10 
a = 8'd95; b = 8'd80;  #10 
a = 8'd95; b = 8'd81;  #10 
a = 8'd95; b = 8'd82;  #10 
a = 8'd95; b = 8'd83;  #10 
a = 8'd95; b = 8'd84;  #10 
a = 8'd95; b = 8'd85;  #10 
a = 8'd95; b = 8'd86;  #10 
a = 8'd95; b = 8'd87;  #10 
a = 8'd95; b = 8'd88;  #10 
a = 8'd95; b = 8'd89;  #10 
a = 8'd95; b = 8'd90;  #10 
a = 8'd95; b = 8'd91;  #10 
a = 8'd95; b = 8'd92;  #10 
a = 8'd95; b = 8'd93;  #10 
a = 8'd95; b = 8'd94;  #10 
a = 8'd95; b = 8'd95;  #10 
a = 8'd95; b = 8'd96;  #10 
a = 8'd95; b = 8'd97;  #10 
a = 8'd95; b = 8'd98;  #10 
a = 8'd95; b = 8'd99;  #10 
a = 8'd95; b = 8'd100;  #10 
a = 8'd95; b = 8'd101;  #10 
a = 8'd95; b = 8'd102;  #10 
a = 8'd95; b = 8'd103;  #10 
a = 8'd95; b = 8'd104;  #10 
a = 8'd95; b = 8'd105;  #10 
a = 8'd95; b = 8'd106;  #10 
a = 8'd95; b = 8'd107;  #10 
a = 8'd95; b = 8'd108;  #10 
a = 8'd95; b = 8'd109;  #10 
a = 8'd95; b = 8'd110;  #10 
a = 8'd95; b = 8'd111;  #10 
a = 8'd95; b = 8'd112;  #10 
a = 8'd95; b = 8'd113;  #10 
a = 8'd95; b = 8'd114;  #10 
a = 8'd95; b = 8'd115;  #10 
a = 8'd95; b = 8'd116;  #10 
a = 8'd95; b = 8'd117;  #10 
a = 8'd95; b = 8'd118;  #10 
a = 8'd95; b = 8'd119;  #10 
a = 8'd95; b = 8'd120;  #10 
a = 8'd95; b = 8'd121;  #10 
a = 8'd95; b = 8'd122;  #10 
a = 8'd95; b = 8'd123;  #10 
a = 8'd95; b = 8'd124;  #10 
a = 8'd95; b = 8'd125;  #10 
a = 8'd95; b = 8'd126;  #10 
a = 8'd95; b = 8'd127;  #10 
a = 8'd95; b = 8'd128;  #10 
a = 8'd95; b = 8'd129;  #10 
a = 8'd95; b = 8'd130;  #10 
a = 8'd95; b = 8'd131;  #10 
a = 8'd95; b = 8'd132;  #10 
a = 8'd95; b = 8'd133;  #10 
a = 8'd95; b = 8'd134;  #10 
a = 8'd95; b = 8'd135;  #10 
a = 8'd95; b = 8'd136;  #10 
a = 8'd95; b = 8'd137;  #10 
a = 8'd95; b = 8'd138;  #10 
a = 8'd95; b = 8'd139;  #10 
a = 8'd95; b = 8'd140;  #10 
a = 8'd95; b = 8'd141;  #10 
a = 8'd95; b = 8'd142;  #10 
a = 8'd95; b = 8'd143;  #10 
a = 8'd95; b = 8'd144;  #10 
a = 8'd95; b = 8'd145;  #10 
a = 8'd95; b = 8'd146;  #10 
a = 8'd95; b = 8'd147;  #10 
a = 8'd95; b = 8'd148;  #10 
a = 8'd95; b = 8'd149;  #10 
a = 8'd95; b = 8'd150;  #10 
a = 8'd95; b = 8'd151;  #10 
a = 8'd95; b = 8'd152;  #10 
a = 8'd95; b = 8'd153;  #10 
a = 8'd95; b = 8'd154;  #10 
a = 8'd95; b = 8'd155;  #10 
a = 8'd95; b = 8'd156;  #10 
a = 8'd95; b = 8'd157;  #10 
a = 8'd95; b = 8'd158;  #10 
a = 8'd95; b = 8'd159;  #10 
a = 8'd95; b = 8'd160;  #10 
a = 8'd95; b = 8'd161;  #10 
a = 8'd95; b = 8'd162;  #10 
a = 8'd95; b = 8'd163;  #10 
a = 8'd95; b = 8'd164;  #10 
a = 8'd95; b = 8'd165;  #10 
a = 8'd95; b = 8'd166;  #10 
a = 8'd95; b = 8'd167;  #10 
a = 8'd95; b = 8'd168;  #10 
a = 8'd95; b = 8'd169;  #10 
a = 8'd95; b = 8'd170;  #10 
a = 8'd95; b = 8'd171;  #10 
a = 8'd95; b = 8'd172;  #10 
a = 8'd95; b = 8'd173;  #10 
a = 8'd95; b = 8'd174;  #10 
a = 8'd95; b = 8'd175;  #10 
a = 8'd95; b = 8'd176;  #10 
a = 8'd95; b = 8'd177;  #10 
a = 8'd95; b = 8'd178;  #10 
a = 8'd95; b = 8'd179;  #10 
a = 8'd95; b = 8'd180;  #10 
a = 8'd95; b = 8'd181;  #10 
a = 8'd95; b = 8'd182;  #10 
a = 8'd95; b = 8'd183;  #10 
a = 8'd95; b = 8'd184;  #10 
a = 8'd95; b = 8'd185;  #10 
a = 8'd95; b = 8'd186;  #10 
a = 8'd95; b = 8'd187;  #10 
a = 8'd95; b = 8'd188;  #10 
a = 8'd95; b = 8'd189;  #10 
a = 8'd95; b = 8'd190;  #10 
a = 8'd95; b = 8'd191;  #10 
a = 8'd95; b = 8'd192;  #10 
a = 8'd95; b = 8'd193;  #10 
a = 8'd95; b = 8'd194;  #10 
a = 8'd95; b = 8'd195;  #10 
a = 8'd95; b = 8'd196;  #10 
a = 8'd95; b = 8'd197;  #10 
a = 8'd95; b = 8'd198;  #10 
a = 8'd95; b = 8'd199;  #10 
a = 8'd95; b = 8'd200;  #10 
a = 8'd95; b = 8'd201;  #10 
a = 8'd95; b = 8'd202;  #10 
a = 8'd95; b = 8'd203;  #10 
a = 8'd95; b = 8'd204;  #10 
a = 8'd95; b = 8'd205;  #10 
a = 8'd95; b = 8'd206;  #10 
a = 8'd95; b = 8'd207;  #10 
a = 8'd95; b = 8'd208;  #10 
a = 8'd95; b = 8'd209;  #10 
a = 8'd95; b = 8'd210;  #10 
a = 8'd95; b = 8'd211;  #10 
a = 8'd95; b = 8'd212;  #10 
a = 8'd95; b = 8'd213;  #10 
a = 8'd95; b = 8'd214;  #10 
a = 8'd95; b = 8'd215;  #10 
a = 8'd95; b = 8'd216;  #10 
a = 8'd95; b = 8'd217;  #10 
a = 8'd95; b = 8'd218;  #10 
a = 8'd95; b = 8'd219;  #10 
a = 8'd95; b = 8'd220;  #10 
a = 8'd95; b = 8'd221;  #10 
a = 8'd95; b = 8'd222;  #10 
a = 8'd95; b = 8'd223;  #10 
a = 8'd95; b = 8'd224;  #10 
a = 8'd95; b = 8'd225;  #10 
a = 8'd95; b = 8'd226;  #10 
a = 8'd95; b = 8'd227;  #10 
a = 8'd95; b = 8'd228;  #10 
a = 8'd95; b = 8'd229;  #10 
a = 8'd95; b = 8'd230;  #10 
a = 8'd95; b = 8'd231;  #10 
a = 8'd95; b = 8'd232;  #10 
a = 8'd95; b = 8'd233;  #10 
a = 8'd95; b = 8'd234;  #10 
a = 8'd95; b = 8'd235;  #10 
a = 8'd95; b = 8'd236;  #10 
a = 8'd95; b = 8'd237;  #10 
a = 8'd95; b = 8'd238;  #10 
a = 8'd95; b = 8'd239;  #10 
a = 8'd95; b = 8'd240;  #10 
a = 8'd95; b = 8'd241;  #10 
a = 8'd95; b = 8'd242;  #10 
a = 8'd95; b = 8'd243;  #10 
a = 8'd95; b = 8'd244;  #10 
a = 8'd95; b = 8'd245;  #10 
a = 8'd95; b = 8'd246;  #10 
a = 8'd95; b = 8'd247;  #10 
a = 8'd95; b = 8'd248;  #10 
a = 8'd95; b = 8'd249;  #10 
a = 8'd95; b = 8'd250;  #10 
a = 8'd95; b = 8'd251;  #10 
a = 8'd95; b = 8'd252;  #10 
a = 8'd95; b = 8'd253;  #10 
a = 8'd95; b = 8'd254;  #10 
a = 8'd95; b = 8'd255;  #10 
a = 8'd96; b = 8'd0;  #10 
a = 8'd96; b = 8'd1;  #10 
a = 8'd96; b = 8'd2;  #10 
a = 8'd96; b = 8'd3;  #10 
a = 8'd96; b = 8'd4;  #10 
a = 8'd96; b = 8'd5;  #10 
a = 8'd96; b = 8'd6;  #10 
a = 8'd96; b = 8'd7;  #10 
a = 8'd96; b = 8'd8;  #10 
a = 8'd96; b = 8'd9;  #10 
a = 8'd96; b = 8'd10;  #10 
a = 8'd96; b = 8'd11;  #10 
a = 8'd96; b = 8'd12;  #10 
a = 8'd96; b = 8'd13;  #10 
a = 8'd96; b = 8'd14;  #10 
a = 8'd96; b = 8'd15;  #10 
a = 8'd96; b = 8'd16;  #10 
a = 8'd96; b = 8'd17;  #10 
a = 8'd96; b = 8'd18;  #10 
a = 8'd96; b = 8'd19;  #10 
a = 8'd96; b = 8'd20;  #10 
a = 8'd96; b = 8'd21;  #10 
a = 8'd96; b = 8'd22;  #10 
a = 8'd96; b = 8'd23;  #10 
a = 8'd96; b = 8'd24;  #10 
a = 8'd96; b = 8'd25;  #10 
a = 8'd96; b = 8'd26;  #10 
a = 8'd96; b = 8'd27;  #10 
a = 8'd96; b = 8'd28;  #10 
a = 8'd96; b = 8'd29;  #10 
a = 8'd96; b = 8'd30;  #10 
a = 8'd96; b = 8'd31;  #10 
a = 8'd96; b = 8'd32;  #10 
a = 8'd96; b = 8'd33;  #10 
a = 8'd96; b = 8'd34;  #10 
a = 8'd96; b = 8'd35;  #10 
a = 8'd96; b = 8'd36;  #10 
a = 8'd96; b = 8'd37;  #10 
a = 8'd96; b = 8'd38;  #10 
a = 8'd96; b = 8'd39;  #10 
a = 8'd96; b = 8'd40;  #10 
a = 8'd96; b = 8'd41;  #10 
a = 8'd96; b = 8'd42;  #10 
a = 8'd96; b = 8'd43;  #10 
a = 8'd96; b = 8'd44;  #10 
a = 8'd96; b = 8'd45;  #10 
a = 8'd96; b = 8'd46;  #10 
a = 8'd96; b = 8'd47;  #10 
a = 8'd96; b = 8'd48;  #10 
a = 8'd96; b = 8'd49;  #10 
a = 8'd96; b = 8'd50;  #10 
a = 8'd96; b = 8'd51;  #10 
a = 8'd96; b = 8'd52;  #10 
a = 8'd96; b = 8'd53;  #10 
a = 8'd96; b = 8'd54;  #10 
a = 8'd96; b = 8'd55;  #10 
a = 8'd96; b = 8'd56;  #10 
a = 8'd96; b = 8'd57;  #10 
a = 8'd96; b = 8'd58;  #10 
a = 8'd96; b = 8'd59;  #10 
a = 8'd96; b = 8'd60;  #10 
a = 8'd96; b = 8'd61;  #10 
a = 8'd96; b = 8'd62;  #10 
a = 8'd96; b = 8'd63;  #10 
a = 8'd96; b = 8'd64;  #10 
a = 8'd96; b = 8'd65;  #10 
a = 8'd96; b = 8'd66;  #10 
a = 8'd96; b = 8'd67;  #10 
a = 8'd96; b = 8'd68;  #10 
a = 8'd96; b = 8'd69;  #10 
a = 8'd96; b = 8'd70;  #10 
a = 8'd96; b = 8'd71;  #10 
a = 8'd96; b = 8'd72;  #10 
a = 8'd96; b = 8'd73;  #10 
a = 8'd96; b = 8'd74;  #10 
a = 8'd96; b = 8'd75;  #10 
a = 8'd96; b = 8'd76;  #10 
a = 8'd96; b = 8'd77;  #10 
a = 8'd96; b = 8'd78;  #10 
a = 8'd96; b = 8'd79;  #10 
a = 8'd96; b = 8'd80;  #10 
a = 8'd96; b = 8'd81;  #10 
a = 8'd96; b = 8'd82;  #10 
a = 8'd96; b = 8'd83;  #10 
a = 8'd96; b = 8'd84;  #10 
a = 8'd96; b = 8'd85;  #10 
a = 8'd96; b = 8'd86;  #10 
a = 8'd96; b = 8'd87;  #10 
a = 8'd96; b = 8'd88;  #10 
a = 8'd96; b = 8'd89;  #10 
a = 8'd96; b = 8'd90;  #10 
a = 8'd96; b = 8'd91;  #10 
a = 8'd96; b = 8'd92;  #10 
a = 8'd96; b = 8'd93;  #10 
a = 8'd96; b = 8'd94;  #10 
a = 8'd96; b = 8'd95;  #10 
a = 8'd96; b = 8'd96;  #10 
a = 8'd96; b = 8'd97;  #10 
a = 8'd96; b = 8'd98;  #10 
a = 8'd96; b = 8'd99;  #10 
a = 8'd96; b = 8'd100;  #10 
a = 8'd96; b = 8'd101;  #10 
a = 8'd96; b = 8'd102;  #10 
a = 8'd96; b = 8'd103;  #10 
a = 8'd96; b = 8'd104;  #10 
a = 8'd96; b = 8'd105;  #10 
a = 8'd96; b = 8'd106;  #10 
a = 8'd96; b = 8'd107;  #10 
a = 8'd96; b = 8'd108;  #10 
a = 8'd96; b = 8'd109;  #10 
a = 8'd96; b = 8'd110;  #10 
a = 8'd96; b = 8'd111;  #10 
a = 8'd96; b = 8'd112;  #10 
a = 8'd96; b = 8'd113;  #10 
a = 8'd96; b = 8'd114;  #10 
a = 8'd96; b = 8'd115;  #10 
a = 8'd96; b = 8'd116;  #10 
a = 8'd96; b = 8'd117;  #10 
a = 8'd96; b = 8'd118;  #10 
a = 8'd96; b = 8'd119;  #10 
a = 8'd96; b = 8'd120;  #10 
a = 8'd96; b = 8'd121;  #10 
a = 8'd96; b = 8'd122;  #10 
a = 8'd96; b = 8'd123;  #10 
a = 8'd96; b = 8'd124;  #10 
a = 8'd96; b = 8'd125;  #10 
a = 8'd96; b = 8'd126;  #10 
a = 8'd96; b = 8'd127;  #10 
a = 8'd96; b = 8'd128;  #10 
a = 8'd96; b = 8'd129;  #10 
a = 8'd96; b = 8'd130;  #10 
a = 8'd96; b = 8'd131;  #10 
a = 8'd96; b = 8'd132;  #10 
a = 8'd96; b = 8'd133;  #10 
a = 8'd96; b = 8'd134;  #10 
a = 8'd96; b = 8'd135;  #10 
a = 8'd96; b = 8'd136;  #10 
a = 8'd96; b = 8'd137;  #10 
a = 8'd96; b = 8'd138;  #10 
a = 8'd96; b = 8'd139;  #10 
a = 8'd96; b = 8'd140;  #10 
a = 8'd96; b = 8'd141;  #10 
a = 8'd96; b = 8'd142;  #10 
a = 8'd96; b = 8'd143;  #10 
a = 8'd96; b = 8'd144;  #10 
a = 8'd96; b = 8'd145;  #10 
a = 8'd96; b = 8'd146;  #10 
a = 8'd96; b = 8'd147;  #10 
a = 8'd96; b = 8'd148;  #10 
a = 8'd96; b = 8'd149;  #10 
a = 8'd96; b = 8'd150;  #10 
a = 8'd96; b = 8'd151;  #10 
a = 8'd96; b = 8'd152;  #10 
a = 8'd96; b = 8'd153;  #10 
a = 8'd96; b = 8'd154;  #10 
a = 8'd96; b = 8'd155;  #10 
a = 8'd96; b = 8'd156;  #10 
a = 8'd96; b = 8'd157;  #10 
a = 8'd96; b = 8'd158;  #10 
a = 8'd96; b = 8'd159;  #10 
a = 8'd96; b = 8'd160;  #10 
a = 8'd96; b = 8'd161;  #10 
a = 8'd96; b = 8'd162;  #10 
a = 8'd96; b = 8'd163;  #10 
a = 8'd96; b = 8'd164;  #10 
a = 8'd96; b = 8'd165;  #10 
a = 8'd96; b = 8'd166;  #10 
a = 8'd96; b = 8'd167;  #10 
a = 8'd96; b = 8'd168;  #10 
a = 8'd96; b = 8'd169;  #10 
a = 8'd96; b = 8'd170;  #10 
a = 8'd96; b = 8'd171;  #10 
a = 8'd96; b = 8'd172;  #10 
a = 8'd96; b = 8'd173;  #10 
a = 8'd96; b = 8'd174;  #10 
a = 8'd96; b = 8'd175;  #10 
a = 8'd96; b = 8'd176;  #10 
a = 8'd96; b = 8'd177;  #10 
a = 8'd96; b = 8'd178;  #10 
a = 8'd96; b = 8'd179;  #10 
a = 8'd96; b = 8'd180;  #10 
a = 8'd96; b = 8'd181;  #10 
a = 8'd96; b = 8'd182;  #10 
a = 8'd96; b = 8'd183;  #10 
a = 8'd96; b = 8'd184;  #10 
a = 8'd96; b = 8'd185;  #10 
a = 8'd96; b = 8'd186;  #10 
a = 8'd96; b = 8'd187;  #10 
a = 8'd96; b = 8'd188;  #10 
a = 8'd96; b = 8'd189;  #10 
a = 8'd96; b = 8'd190;  #10 
a = 8'd96; b = 8'd191;  #10 
a = 8'd96; b = 8'd192;  #10 
a = 8'd96; b = 8'd193;  #10 
a = 8'd96; b = 8'd194;  #10 
a = 8'd96; b = 8'd195;  #10 
a = 8'd96; b = 8'd196;  #10 
a = 8'd96; b = 8'd197;  #10 
a = 8'd96; b = 8'd198;  #10 
a = 8'd96; b = 8'd199;  #10 
a = 8'd96; b = 8'd200;  #10 
a = 8'd96; b = 8'd201;  #10 
a = 8'd96; b = 8'd202;  #10 
a = 8'd96; b = 8'd203;  #10 
a = 8'd96; b = 8'd204;  #10 
a = 8'd96; b = 8'd205;  #10 
a = 8'd96; b = 8'd206;  #10 
a = 8'd96; b = 8'd207;  #10 
a = 8'd96; b = 8'd208;  #10 
a = 8'd96; b = 8'd209;  #10 
a = 8'd96; b = 8'd210;  #10 
a = 8'd96; b = 8'd211;  #10 
a = 8'd96; b = 8'd212;  #10 
a = 8'd96; b = 8'd213;  #10 
a = 8'd96; b = 8'd214;  #10 
a = 8'd96; b = 8'd215;  #10 
a = 8'd96; b = 8'd216;  #10 
a = 8'd96; b = 8'd217;  #10 
a = 8'd96; b = 8'd218;  #10 
a = 8'd96; b = 8'd219;  #10 
a = 8'd96; b = 8'd220;  #10 
a = 8'd96; b = 8'd221;  #10 
a = 8'd96; b = 8'd222;  #10 
a = 8'd96; b = 8'd223;  #10 
a = 8'd96; b = 8'd224;  #10 
a = 8'd96; b = 8'd225;  #10 
a = 8'd96; b = 8'd226;  #10 
a = 8'd96; b = 8'd227;  #10 
a = 8'd96; b = 8'd228;  #10 
a = 8'd96; b = 8'd229;  #10 
a = 8'd96; b = 8'd230;  #10 
a = 8'd96; b = 8'd231;  #10 
a = 8'd96; b = 8'd232;  #10 
a = 8'd96; b = 8'd233;  #10 
a = 8'd96; b = 8'd234;  #10 
a = 8'd96; b = 8'd235;  #10 
a = 8'd96; b = 8'd236;  #10 
a = 8'd96; b = 8'd237;  #10 
a = 8'd96; b = 8'd238;  #10 
a = 8'd96; b = 8'd239;  #10 
a = 8'd96; b = 8'd240;  #10 
a = 8'd96; b = 8'd241;  #10 
a = 8'd96; b = 8'd242;  #10 
a = 8'd96; b = 8'd243;  #10 
a = 8'd96; b = 8'd244;  #10 
a = 8'd96; b = 8'd245;  #10 
a = 8'd96; b = 8'd246;  #10 
a = 8'd96; b = 8'd247;  #10 
a = 8'd96; b = 8'd248;  #10 
a = 8'd96; b = 8'd249;  #10 
a = 8'd96; b = 8'd250;  #10 
a = 8'd96; b = 8'd251;  #10 
a = 8'd96; b = 8'd252;  #10 
a = 8'd96; b = 8'd253;  #10 
a = 8'd96; b = 8'd254;  #10 
a = 8'd96; b = 8'd255;  #10 
a = 8'd97; b = 8'd0;  #10 
a = 8'd97; b = 8'd1;  #10 
a = 8'd97; b = 8'd2;  #10 
a = 8'd97; b = 8'd3;  #10 
a = 8'd97; b = 8'd4;  #10 
a = 8'd97; b = 8'd5;  #10 
a = 8'd97; b = 8'd6;  #10 
a = 8'd97; b = 8'd7;  #10 
a = 8'd97; b = 8'd8;  #10 
a = 8'd97; b = 8'd9;  #10 
a = 8'd97; b = 8'd10;  #10 
a = 8'd97; b = 8'd11;  #10 
a = 8'd97; b = 8'd12;  #10 
a = 8'd97; b = 8'd13;  #10 
a = 8'd97; b = 8'd14;  #10 
a = 8'd97; b = 8'd15;  #10 
a = 8'd97; b = 8'd16;  #10 
a = 8'd97; b = 8'd17;  #10 
a = 8'd97; b = 8'd18;  #10 
a = 8'd97; b = 8'd19;  #10 
a = 8'd97; b = 8'd20;  #10 
a = 8'd97; b = 8'd21;  #10 
a = 8'd97; b = 8'd22;  #10 
a = 8'd97; b = 8'd23;  #10 
a = 8'd97; b = 8'd24;  #10 
a = 8'd97; b = 8'd25;  #10 
a = 8'd97; b = 8'd26;  #10 
a = 8'd97; b = 8'd27;  #10 
a = 8'd97; b = 8'd28;  #10 
a = 8'd97; b = 8'd29;  #10 
a = 8'd97; b = 8'd30;  #10 
a = 8'd97; b = 8'd31;  #10 
a = 8'd97; b = 8'd32;  #10 
a = 8'd97; b = 8'd33;  #10 
a = 8'd97; b = 8'd34;  #10 
a = 8'd97; b = 8'd35;  #10 
a = 8'd97; b = 8'd36;  #10 
a = 8'd97; b = 8'd37;  #10 
a = 8'd97; b = 8'd38;  #10 
a = 8'd97; b = 8'd39;  #10 
a = 8'd97; b = 8'd40;  #10 
a = 8'd97; b = 8'd41;  #10 
a = 8'd97; b = 8'd42;  #10 
a = 8'd97; b = 8'd43;  #10 
a = 8'd97; b = 8'd44;  #10 
a = 8'd97; b = 8'd45;  #10 
a = 8'd97; b = 8'd46;  #10 
a = 8'd97; b = 8'd47;  #10 
a = 8'd97; b = 8'd48;  #10 
a = 8'd97; b = 8'd49;  #10 
a = 8'd97; b = 8'd50;  #10 
a = 8'd97; b = 8'd51;  #10 
a = 8'd97; b = 8'd52;  #10 
a = 8'd97; b = 8'd53;  #10 
a = 8'd97; b = 8'd54;  #10 
a = 8'd97; b = 8'd55;  #10 
a = 8'd97; b = 8'd56;  #10 
a = 8'd97; b = 8'd57;  #10 
a = 8'd97; b = 8'd58;  #10 
a = 8'd97; b = 8'd59;  #10 
a = 8'd97; b = 8'd60;  #10 
a = 8'd97; b = 8'd61;  #10 
a = 8'd97; b = 8'd62;  #10 
a = 8'd97; b = 8'd63;  #10 
a = 8'd97; b = 8'd64;  #10 
a = 8'd97; b = 8'd65;  #10 
a = 8'd97; b = 8'd66;  #10 
a = 8'd97; b = 8'd67;  #10 
a = 8'd97; b = 8'd68;  #10 
a = 8'd97; b = 8'd69;  #10 
a = 8'd97; b = 8'd70;  #10 
a = 8'd97; b = 8'd71;  #10 
a = 8'd97; b = 8'd72;  #10 
a = 8'd97; b = 8'd73;  #10 
a = 8'd97; b = 8'd74;  #10 
a = 8'd97; b = 8'd75;  #10 
a = 8'd97; b = 8'd76;  #10 
a = 8'd97; b = 8'd77;  #10 
a = 8'd97; b = 8'd78;  #10 
a = 8'd97; b = 8'd79;  #10 
a = 8'd97; b = 8'd80;  #10 
a = 8'd97; b = 8'd81;  #10 
a = 8'd97; b = 8'd82;  #10 
a = 8'd97; b = 8'd83;  #10 
a = 8'd97; b = 8'd84;  #10 
a = 8'd97; b = 8'd85;  #10 
a = 8'd97; b = 8'd86;  #10 
a = 8'd97; b = 8'd87;  #10 
a = 8'd97; b = 8'd88;  #10 
a = 8'd97; b = 8'd89;  #10 
a = 8'd97; b = 8'd90;  #10 
a = 8'd97; b = 8'd91;  #10 
a = 8'd97; b = 8'd92;  #10 
a = 8'd97; b = 8'd93;  #10 
a = 8'd97; b = 8'd94;  #10 
a = 8'd97; b = 8'd95;  #10 
a = 8'd97; b = 8'd96;  #10 
a = 8'd97; b = 8'd97;  #10 
a = 8'd97; b = 8'd98;  #10 
a = 8'd97; b = 8'd99;  #10 
a = 8'd97; b = 8'd100;  #10 
a = 8'd97; b = 8'd101;  #10 
a = 8'd97; b = 8'd102;  #10 
a = 8'd97; b = 8'd103;  #10 
a = 8'd97; b = 8'd104;  #10 
a = 8'd97; b = 8'd105;  #10 
a = 8'd97; b = 8'd106;  #10 
a = 8'd97; b = 8'd107;  #10 
a = 8'd97; b = 8'd108;  #10 
a = 8'd97; b = 8'd109;  #10 
a = 8'd97; b = 8'd110;  #10 
a = 8'd97; b = 8'd111;  #10 
a = 8'd97; b = 8'd112;  #10 
a = 8'd97; b = 8'd113;  #10 
a = 8'd97; b = 8'd114;  #10 
a = 8'd97; b = 8'd115;  #10 
a = 8'd97; b = 8'd116;  #10 
a = 8'd97; b = 8'd117;  #10 
a = 8'd97; b = 8'd118;  #10 
a = 8'd97; b = 8'd119;  #10 
a = 8'd97; b = 8'd120;  #10 
a = 8'd97; b = 8'd121;  #10 
a = 8'd97; b = 8'd122;  #10 
a = 8'd97; b = 8'd123;  #10 
a = 8'd97; b = 8'd124;  #10 
a = 8'd97; b = 8'd125;  #10 
a = 8'd97; b = 8'd126;  #10 
a = 8'd97; b = 8'd127;  #10 
a = 8'd97; b = 8'd128;  #10 
a = 8'd97; b = 8'd129;  #10 
a = 8'd97; b = 8'd130;  #10 
a = 8'd97; b = 8'd131;  #10 
a = 8'd97; b = 8'd132;  #10 
a = 8'd97; b = 8'd133;  #10 
a = 8'd97; b = 8'd134;  #10 
a = 8'd97; b = 8'd135;  #10 
a = 8'd97; b = 8'd136;  #10 
a = 8'd97; b = 8'd137;  #10 
a = 8'd97; b = 8'd138;  #10 
a = 8'd97; b = 8'd139;  #10 
a = 8'd97; b = 8'd140;  #10 
a = 8'd97; b = 8'd141;  #10 
a = 8'd97; b = 8'd142;  #10 
a = 8'd97; b = 8'd143;  #10 
a = 8'd97; b = 8'd144;  #10 
a = 8'd97; b = 8'd145;  #10 
a = 8'd97; b = 8'd146;  #10 
a = 8'd97; b = 8'd147;  #10 
a = 8'd97; b = 8'd148;  #10 
a = 8'd97; b = 8'd149;  #10 
a = 8'd97; b = 8'd150;  #10 
a = 8'd97; b = 8'd151;  #10 
a = 8'd97; b = 8'd152;  #10 
a = 8'd97; b = 8'd153;  #10 
a = 8'd97; b = 8'd154;  #10 
a = 8'd97; b = 8'd155;  #10 
a = 8'd97; b = 8'd156;  #10 
a = 8'd97; b = 8'd157;  #10 
a = 8'd97; b = 8'd158;  #10 
a = 8'd97; b = 8'd159;  #10 
a = 8'd97; b = 8'd160;  #10 
a = 8'd97; b = 8'd161;  #10 
a = 8'd97; b = 8'd162;  #10 
a = 8'd97; b = 8'd163;  #10 
a = 8'd97; b = 8'd164;  #10 
a = 8'd97; b = 8'd165;  #10 
a = 8'd97; b = 8'd166;  #10 
a = 8'd97; b = 8'd167;  #10 
a = 8'd97; b = 8'd168;  #10 
a = 8'd97; b = 8'd169;  #10 
a = 8'd97; b = 8'd170;  #10 
a = 8'd97; b = 8'd171;  #10 
a = 8'd97; b = 8'd172;  #10 
a = 8'd97; b = 8'd173;  #10 
a = 8'd97; b = 8'd174;  #10 
a = 8'd97; b = 8'd175;  #10 
a = 8'd97; b = 8'd176;  #10 
a = 8'd97; b = 8'd177;  #10 
a = 8'd97; b = 8'd178;  #10 
a = 8'd97; b = 8'd179;  #10 
a = 8'd97; b = 8'd180;  #10 
a = 8'd97; b = 8'd181;  #10 
a = 8'd97; b = 8'd182;  #10 
a = 8'd97; b = 8'd183;  #10 
a = 8'd97; b = 8'd184;  #10 
a = 8'd97; b = 8'd185;  #10 
a = 8'd97; b = 8'd186;  #10 
a = 8'd97; b = 8'd187;  #10 
a = 8'd97; b = 8'd188;  #10 
a = 8'd97; b = 8'd189;  #10 
a = 8'd97; b = 8'd190;  #10 
a = 8'd97; b = 8'd191;  #10 
a = 8'd97; b = 8'd192;  #10 
a = 8'd97; b = 8'd193;  #10 
a = 8'd97; b = 8'd194;  #10 
a = 8'd97; b = 8'd195;  #10 
a = 8'd97; b = 8'd196;  #10 
a = 8'd97; b = 8'd197;  #10 
a = 8'd97; b = 8'd198;  #10 
a = 8'd97; b = 8'd199;  #10 
a = 8'd97; b = 8'd200;  #10 
a = 8'd97; b = 8'd201;  #10 
a = 8'd97; b = 8'd202;  #10 
a = 8'd97; b = 8'd203;  #10 
a = 8'd97; b = 8'd204;  #10 
a = 8'd97; b = 8'd205;  #10 
a = 8'd97; b = 8'd206;  #10 
a = 8'd97; b = 8'd207;  #10 
a = 8'd97; b = 8'd208;  #10 
a = 8'd97; b = 8'd209;  #10 
a = 8'd97; b = 8'd210;  #10 
a = 8'd97; b = 8'd211;  #10 
a = 8'd97; b = 8'd212;  #10 
a = 8'd97; b = 8'd213;  #10 
a = 8'd97; b = 8'd214;  #10 
a = 8'd97; b = 8'd215;  #10 
a = 8'd97; b = 8'd216;  #10 
a = 8'd97; b = 8'd217;  #10 
a = 8'd97; b = 8'd218;  #10 
a = 8'd97; b = 8'd219;  #10 
a = 8'd97; b = 8'd220;  #10 
a = 8'd97; b = 8'd221;  #10 
a = 8'd97; b = 8'd222;  #10 
a = 8'd97; b = 8'd223;  #10 
a = 8'd97; b = 8'd224;  #10 
a = 8'd97; b = 8'd225;  #10 
a = 8'd97; b = 8'd226;  #10 
a = 8'd97; b = 8'd227;  #10 
a = 8'd97; b = 8'd228;  #10 
a = 8'd97; b = 8'd229;  #10 
a = 8'd97; b = 8'd230;  #10 
a = 8'd97; b = 8'd231;  #10 
a = 8'd97; b = 8'd232;  #10 
a = 8'd97; b = 8'd233;  #10 
a = 8'd97; b = 8'd234;  #10 
a = 8'd97; b = 8'd235;  #10 
a = 8'd97; b = 8'd236;  #10 
a = 8'd97; b = 8'd237;  #10 
a = 8'd97; b = 8'd238;  #10 
a = 8'd97; b = 8'd239;  #10 
a = 8'd97; b = 8'd240;  #10 
a = 8'd97; b = 8'd241;  #10 
a = 8'd97; b = 8'd242;  #10 
a = 8'd97; b = 8'd243;  #10 
a = 8'd97; b = 8'd244;  #10 
a = 8'd97; b = 8'd245;  #10 
a = 8'd97; b = 8'd246;  #10 
a = 8'd97; b = 8'd247;  #10 
a = 8'd97; b = 8'd248;  #10 
a = 8'd97; b = 8'd249;  #10 
a = 8'd97; b = 8'd250;  #10 
a = 8'd97; b = 8'd251;  #10 
a = 8'd97; b = 8'd252;  #10 
a = 8'd97; b = 8'd253;  #10 
a = 8'd97; b = 8'd254;  #10 
a = 8'd97; b = 8'd255;  #10 
a = 8'd98; b = 8'd0;  #10 
a = 8'd98; b = 8'd1;  #10 
a = 8'd98; b = 8'd2;  #10 
a = 8'd98; b = 8'd3;  #10 
a = 8'd98; b = 8'd4;  #10 
a = 8'd98; b = 8'd5;  #10 
a = 8'd98; b = 8'd6;  #10 
a = 8'd98; b = 8'd7;  #10 
a = 8'd98; b = 8'd8;  #10 
a = 8'd98; b = 8'd9;  #10 
a = 8'd98; b = 8'd10;  #10 
a = 8'd98; b = 8'd11;  #10 
a = 8'd98; b = 8'd12;  #10 
a = 8'd98; b = 8'd13;  #10 
a = 8'd98; b = 8'd14;  #10 
a = 8'd98; b = 8'd15;  #10 
a = 8'd98; b = 8'd16;  #10 
a = 8'd98; b = 8'd17;  #10 
a = 8'd98; b = 8'd18;  #10 
a = 8'd98; b = 8'd19;  #10 
a = 8'd98; b = 8'd20;  #10 
a = 8'd98; b = 8'd21;  #10 
a = 8'd98; b = 8'd22;  #10 
a = 8'd98; b = 8'd23;  #10 
a = 8'd98; b = 8'd24;  #10 
a = 8'd98; b = 8'd25;  #10 
a = 8'd98; b = 8'd26;  #10 
a = 8'd98; b = 8'd27;  #10 
a = 8'd98; b = 8'd28;  #10 
a = 8'd98; b = 8'd29;  #10 
a = 8'd98; b = 8'd30;  #10 
a = 8'd98; b = 8'd31;  #10 
a = 8'd98; b = 8'd32;  #10 
a = 8'd98; b = 8'd33;  #10 
a = 8'd98; b = 8'd34;  #10 
a = 8'd98; b = 8'd35;  #10 
a = 8'd98; b = 8'd36;  #10 
a = 8'd98; b = 8'd37;  #10 
a = 8'd98; b = 8'd38;  #10 
a = 8'd98; b = 8'd39;  #10 
a = 8'd98; b = 8'd40;  #10 
a = 8'd98; b = 8'd41;  #10 
a = 8'd98; b = 8'd42;  #10 
a = 8'd98; b = 8'd43;  #10 
a = 8'd98; b = 8'd44;  #10 
a = 8'd98; b = 8'd45;  #10 
a = 8'd98; b = 8'd46;  #10 
a = 8'd98; b = 8'd47;  #10 
a = 8'd98; b = 8'd48;  #10 
a = 8'd98; b = 8'd49;  #10 
a = 8'd98; b = 8'd50;  #10 
a = 8'd98; b = 8'd51;  #10 
a = 8'd98; b = 8'd52;  #10 
a = 8'd98; b = 8'd53;  #10 
a = 8'd98; b = 8'd54;  #10 
a = 8'd98; b = 8'd55;  #10 
a = 8'd98; b = 8'd56;  #10 
a = 8'd98; b = 8'd57;  #10 
a = 8'd98; b = 8'd58;  #10 
a = 8'd98; b = 8'd59;  #10 
a = 8'd98; b = 8'd60;  #10 
a = 8'd98; b = 8'd61;  #10 
a = 8'd98; b = 8'd62;  #10 
a = 8'd98; b = 8'd63;  #10 
a = 8'd98; b = 8'd64;  #10 
a = 8'd98; b = 8'd65;  #10 
a = 8'd98; b = 8'd66;  #10 
a = 8'd98; b = 8'd67;  #10 
a = 8'd98; b = 8'd68;  #10 
a = 8'd98; b = 8'd69;  #10 
a = 8'd98; b = 8'd70;  #10 
a = 8'd98; b = 8'd71;  #10 
a = 8'd98; b = 8'd72;  #10 
a = 8'd98; b = 8'd73;  #10 
a = 8'd98; b = 8'd74;  #10 
a = 8'd98; b = 8'd75;  #10 
a = 8'd98; b = 8'd76;  #10 
a = 8'd98; b = 8'd77;  #10 
a = 8'd98; b = 8'd78;  #10 
a = 8'd98; b = 8'd79;  #10 
a = 8'd98; b = 8'd80;  #10 
a = 8'd98; b = 8'd81;  #10 
a = 8'd98; b = 8'd82;  #10 
a = 8'd98; b = 8'd83;  #10 
a = 8'd98; b = 8'd84;  #10 
a = 8'd98; b = 8'd85;  #10 
a = 8'd98; b = 8'd86;  #10 
a = 8'd98; b = 8'd87;  #10 
a = 8'd98; b = 8'd88;  #10 
a = 8'd98; b = 8'd89;  #10 
a = 8'd98; b = 8'd90;  #10 
a = 8'd98; b = 8'd91;  #10 
a = 8'd98; b = 8'd92;  #10 
a = 8'd98; b = 8'd93;  #10 
a = 8'd98; b = 8'd94;  #10 
a = 8'd98; b = 8'd95;  #10 
a = 8'd98; b = 8'd96;  #10 
a = 8'd98; b = 8'd97;  #10 
a = 8'd98; b = 8'd98;  #10 
a = 8'd98; b = 8'd99;  #10 
a = 8'd98; b = 8'd100;  #10 
a = 8'd98; b = 8'd101;  #10 
a = 8'd98; b = 8'd102;  #10 
a = 8'd98; b = 8'd103;  #10 
a = 8'd98; b = 8'd104;  #10 
a = 8'd98; b = 8'd105;  #10 
a = 8'd98; b = 8'd106;  #10 
a = 8'd98; b = 8'd107;  #10 
a = 8'd98; b = 8'd108;  #10 
a = 8'd98; b = 8'd109;  #10 
a = 8'd98; b = 8'd110;  #10 
a = 8'd98; b = 8'd111;  #10 
a = 8'd98; b = 8'd112;  #10 
a = 8'd98; b = 8'd113;  #10 
a = 8'd98; b = 8'd114;  #10 
a = 8'd98; b = 8'd115;  #10 
a = 8'd98; b = 8'd116;  #10 
a = 8'd98; b = 8'd117;  #10 
a = 8'd98; b = 8'd118;  #10 
a = 8'd98; b = 8'd119;  #10 
a = 8'd98; b = 8'd120;  #10 
a = 8'd98; b = 8'd121;  #10 
a = 8'd98; b = 8'd122;  #10 
a = 8'd98; b = 8'd123;  #10 
a = 8'd98; b = 8'd124;  #10 
a = 8'd98; b = 8'd125;  #10 
a = 8'd98; b = 8'd126;  #10 
a = 8'd98; b = 8'd127;  #10 
a = 8'd98; b = 8'd128;  #10 
a = 8'd98; b = 8'd129;  #10 
a = 8'd98; b = 8'd130;  #10 
a = 8'd98; b = 8'd131;  #10 
a = 8'd98; b = 8'd132;  #10 
a = 8'd98; b = 8'd133;  #10 
a = 8'd98; b = 8'd134;  #10 
a = 8'd98; b = 8'd135;  #10 
a = 8'd98; b = 8'd136;  #10 
a = 8'd98; b = 8'd137;  #10 
a = 8'd98; b = 8'd138;  #10 
a = 8'd98; b = 8'd139;  #10 
a = 8'd98; b = 8'd140;  #10 
a = 8'd98; b = 8'd141;  #10 
a = 8'd98; b = 8'd142;  #10 
a = 8'd98; b = 8'd143;  #10 
a = 8'd98; b = 8'd144;  #10 
a = 8'd98; b = 8'd145;  #10 
a = 8'd98; b = 8'd146;  #10 
a = 8'd98; b = 8'd147;  #10 
a = 8'd98; b = 8'd148;  #10 
a = 8'd98; b = 8'd149;  #10 
a = 8'd98; b = 8'd150;  #10 
a = 8'd98; b = 8'd151;  #10 
a = 8'd98; b = 8'd152;  #10 
a = 8'd98; b = 8'd153;  #10 
a = 8'd98; b = 8'd154;  #10 
a = 8'd98; b = 8'd155;  #10 
a = 8'd98; b = 8'd156;  #10 
a = 8'd98; b = 8'd157;  #10 
a = 8'd98; b = 8'd158;  #10 
a = 8'd98; b = 8'd159;  #10 
a = 8'd98; b = 8'd160;  #10 
a = 8'd98; b = 8'd161;  #10 
a = 8'd98; b = 8'd162;  #10 
a = 8'd98; b = 8'd163;  #10 
a = 8'd98; b = 8'd164;  #10 
a = 8'd98; b = 8'd165;  #10 
a = 8'd98; b = 8'd166;  #10 
a = 8'd98; b = 8'd167;  #10 
a = 8'd98; b = 8'd168;  #10 
a = 8'd98; b = 8'd169;  #10 
a = 8'd98; b = 8'd170;  #10 
a = 8'd98; b = 8'd171;  #10 
a = 8'd98; b = 8'd172;  #10 
a = 8'd98; b = 8'd173;  #10 
a = 8'd98; b = 8'd174;  #10 
a = 8'd98; b = 8'd175;  #10 
a = 8'd98; b = 8'd176;  #10 
a = 8'd98; b = 8'd177;  #10 
a = 8'd98; b = 8'd178;  #10 
a = 8'd98; b = 8'd179;  #10 
a = 8'd98; b = 8'd180;  #10 
a = 8'd98; b = 8'd181;  #10 
a = 8'd98; b = 8'd182;  #10 
a = 8'd98; b = 8'd183;  #10 
a = 8'd98; b = 8'd184;  #10 
a = 8'd98; b = 8'd185;  #10 
a = 8'd98; b = 8'd186;  #10 
a = 8'd98; b = 8'd187;  #10 
a = 8'd98; b = 8'd188;  #10 
a = 8'd98; b = 8'd189;  #10 
a = 8'd98; b = 8'd190;  #10 
a = 8'd98; b = 8'd191;  #10 
a = 8'd98; b = 8'd192;  #10 
a = 8'd98; b = 8'd193;  #10 
a = 8'd98; b = 8'd194;  #10 
a = 8'd98; b = 8'd195;  #10 
a = 8'd98; b = 8'd196;  #10 
a = 8'd98; b = 8'd197;  #10 
a = 8'd98; b = 8'd198;  #10 
a = 8'd98; b = 8'd199;  #10 
a = 8'd98; b = 8'd200;  #10 
a = 8'd98; b = 8'd201;  #10 
a = 8'd98; b = 8'd202;  #10 
a = 8'd98; b = 8'd203;  #10 
a = 8'd98; b = 8'd204;  #10 
a = 8'd98; b = 8'd205;  #10 
a = 8'd98; b = 8'd206;  #10 
a = 8'd98; b = 8'd207;  #10 
a = 8'd98; b = 8'd208;  #10 
a = 8'd98; b = 8'd209;  #10 
a = 8'd98; b = 8'd210;  #10 
a = 8'd98; b = 8'd211;  #10 
a = 8'd98; b = 8'd212;  #10 
a = 8'd98; b = 8'd213;  #10 
a = 8'd98; b = 8'd214;  #10 
a = 8'd98; b = 8'd215;  #10 
a = 8'd98; b = 8'd216;  #10 
a = 8'd98; b = 8'd217;  #10 
a = 8'd98; b = 8'd218;  #10 
a = 8'd98; b = 8'd219;  #10 
a = 8'd98; b = 8'd220;  #10 
a = 8'd98; b = 8'd221;  #10 
a = 8'd98; b = 8'd222;  #10 
a = 8'd98; b = 8'd223;  #10 
a = 8'd98; b = 8'd224;  #10 
a = 8'd98; b = 8'd225;  #10 
a = 8'd98; b = 8'd226;  #10 
a = 8'd98; b = 8'd227;  #10 
a = 8'd98; b = 8'd228;  #10 
a = 8'd98; b = 8'd229;  #10 
a = 8'd98; b = 8'd230;  #10 
a = 8'd98; b = 8'd231;  #10 
a = 8'd98; b = 8'd232;  #10 
a = 8'd98; b = 8'd233;  #10 
a = 8'd98; b = 8'd234;  #10 
a = 8'd98; b = 8'd235;  #10 
a = 8'd98; b = 8'd236;  #10 
a = 8'd98; b = 8'd237;  #10 
a = 8'd98; b = 8'd238;  #10 
a = 8'd98; b = 8'd239;  #10 
a = 8'd98; b = 8'd240;  #10 
a = 8'd98; b = 8'd241;  #10 
a = 8'd98; b = 8'd242;  #10 
a = 8'd98; b = 8'd243;  #10 
a = 8'd98; b = 8'd244;  #10 
a = 8'd98; b = 8'd245;  #10 
a = 8'd98; b = 8'd246;  #10 
a = 8'd98; b = 8'd247;  #10 
a = 8'd98; b = 8'd248;  #10 
a = 8'd98; b = 8'd249;  #10 
a = 8'd98; b = 8'd250;  #10 
a = 8'd98; b = 8'd251;  #10 
a = 8'd98; b = 8'd252;  #10 
a = 8'd98; b = 8'd253;  #10 
a = 8'd98; b = 8'd254;  #10 
a = 8'd98; b = 8'd255;  #10 
a = 8'd99; b = 8'd0;  #10 
a = 8'd99; b = 8'd1;  #10 
a = 8'd99; b = 8'd2;  #10 
a = 8'd99; b = 8'd3;  #10 
a = 8'd99; b = 8'd4;  #10 
a = 8'd99; b = 8'd5;  #10 
a = 8'd99; b = 8'd6;  #10 
a = 8'd99; b = 8'd7;  #10 
a = 8'd99; b = 8'd8;  #10 
a = 8'd99; b = 8'd9;  #10 
a = 8'd99; b = 8'd10;  #10 
a = 8'd99; b = 8'd11;  #10 
a = 8'd99; b = 8'd12;  #10 
a = 8'd99; b = 8'd13;  #10 
a = 8'd99; b = 8'd14;  #10 
a = 8'd99; b = 8'd15;  #10 
a = 8'd99; b = 8'd16;  #10 
a = 8'd99; b = 8'd17;  #10 
a = 8'd99; b = 8'd18;  #10 
a = 8'd99; b = 8'd19;  #10 
a = 8'd99; b = 8'd20;  #10 
a = 8'd99; b = 8'd21;  #10 
a = 8'd99; b = 8'd22;  #10 
a = 8'd99; b = 8'd23;  #10 
a = 8'd99; b = 8'd24;  #10 
a = 8'd99; b = 8'd25;  #10 
a = 8'd99; b = 8'd26;  #10 
a = 8'd99; b = 8'd27;  #10 
a = 8'd99; b = 8'd28;  #10 
a = 8'd99; b = 8'd29;  #10 
a = 8'd99; b = 8'd30;  #10 
a = 8'd99; b = 8'd31;  #10 
a = 8'd99; b = 8'd32;  #10 
a = 8'd99; b = 8'd33;  #10 
a = 8'd99; b = 8'd34;  #10 
a = 8'd99; b = 8'd35;  #10 
a = 8'd99; b = 8'd36;  #10 
a = 8'd99; b = 8'd37;  #10 
a = 8'd99; b = 8'd38;  #10 
a = 8'd99; b = 8'd39;  #10 
a = 8'd99; b = 8'd40;  #10 
a = 8'd99; b = 8'd41;  #10 
a = 8'd99; b = 8'd42;  #10 
a = 8'd99; b = 8'd43;  #10 
a = 8'd99; b = 8'd44;  #10 
a = 8'd99; b = 8'd45;  #10 
a = 8'd99; b = 8'd46;  #10 
a = 8'd99; b = 8'd47;  #10 
a = 8'd99; b = 8'd48;  #10 
a = 8'd99; b = 8'd49;  #10 
a = 8'd99; b = 8'd50;  #10 
a = 8'd99; b = 8'd51;  #10 
a = 8'd99; b = 8'd52;  #10 
a = 8'd99; b = 8'd53;  #10 
a = 8'd99; b = 8'd54;  #10 
a = 8'd99; b = 8'd55;  #10 
a = 8'd99; b = 8'd56;  #10 
a = 8'd99; b = 8'd57;  #10 
a = 8'd99; b = 8'd58;  #10 
a = 8'd99; b = 8'd59;  #10 
a = 8'd99; b = 8'd60;  #10 
a = 8'd99; b = 8'd61;  #10 
a = 8'd99; b = 8'd62;  #10 
a = 8'd99; b = 8'd63;  #10 
a = 8'd99; b = 8'd64;  #10 
a = 8'd99; b = 8'd65;  #10 
a = 8'd99; b = 8'd66;  #10 
a = 8'd99; b = 8'd67;  #10 
a = 8'd99; b = 8'd68;  #10 
a = 8'd99; b = 8'd69;  #10 
a = 8'd99; b = 8'd70;  #10 
a = 8'd99; b = 8'd71;  #10 
a = 8'd99; b = 8'd72;  #10 
a = 8'd99; b = 8'd73;  #10 
a = 8'd99; b = 8'd74;  #10 
a = 8'd99; b = 8'd75;  #10 
a = 8'd99; b = 8'd76;  #10 
a = 8'd99; b = 8'd77;  #10 
a = 8'd99; b = 8'd78;  #10 
a = 8'd99; b = 8'd79;  #10 
a = 8'd99; b = 8'd80;  #10 
a = 8'd99; b = 8'd81;  #10 
a = 8'd99; b = 8'd82;  #10 
a = 8'd99; b = 8'd83;  #10 
a = 8'd99; b = 8'd84;  #10 
a = 8'd99; b = 8'd85;  #10 
a = 8'd99; b = 8'd86;  #10 
a = 8'd99; b = 8'd87;  #10 
a = 8'd99; b = 8'd88;  #10 
a = 8'd99; b = 8'd89;  #10 
a = 8'd99; b = 8'd90;  #10 
a = 8'd99; b = 8'd91;  #10 
a = 8'd99; b = 8'd92;  #10 
a = 8'd99; b = 8'd93;  #10 
a = 8'd99; b = 8'd94;  #10 
a = 8'd99; b = 8'd95;  #10 
a = 8'd99; b = 8'd96;  #10 
a = 8'd99; b = 8'd97;  #10 
a = 8'd99; b = 8'd98;  #10 
a = 8'd99; b = 8'd99;  #10 
a = 8'd99; b = 8'd100;  #10 
a = 8'd99; b = 8'd101;  #10 
a = 8'd99; b = 8'd102;  #10 
a = 8'd99; b = 8'd103;  #10 
a = 8'd99; b = 8'd104;  #10 
a = 8'd99; b = 8'd105;  #10 
a = 8'd99; b = 8'd106;  #10 
a = 8'd99; b = 8'd107;  #10 
a = 8'd99; b = 8'd108;  #10 
a = 8'd99; b = 8'd109;  #10 
a = 8'd99; b = 8'd110;  #10 
a = 8'd99; b = 8'd111;  #10 
a = 8'd99; b = 8'd112;  #10 
a = 8'd99; b = 8'd113;  #10 
a = 8'd99; b = 8'd114;  #10 
a = 8'd99; b = 8'd115;  #10 
a = 8'd99; b = 8'd116;  #10 
a = 8'd99; b = 8'd117;  #10 
a = 8'd99; b = 8'd118;  #10 
a = 8'd99; b = 8'd119;  #10 
a = 8'd99; b = 8'd120;  #10 
a = 8'd99; b = 8'd121;  #10 
a = 8'd99; b = 8'd122;  #10 
a = 8'd99; b = 8'd123;  #10 
a = 8'd99; b = 8'd124;  #10 
a = 8'd99; b = 8'd125;  #10 
a = 8'd99; b = 8'd126;  #10 
a = 8'd99; b = 8'd127;  #10 
a = 8'd99; b = 8'd128;  #10 
a = 8'd99; b = 8'd129;  #10 
a = 8'd99; b = 8'd130;  #10 
a = 8'd99; b = 8'd131;  #10 
a = 8'd99; b = 8'd132;  #10 
a = 8'd99; b = 8'd133;  #10 
a = 8'd99; b = 8'd134;  #10 
a = 8'd99; b = 8'd135;  #10 
a = 8'd99; b = 8'd136;  #10 
a = 8'd99; b = 8'd137;  #10 
a = 8'd99; b = 8'd138;  #10 
a = 8'd99; b = 8'd139;  #10 
a = 8'd99; b = 8'd140;  #10 
a = 8'd99; b = 8'd141;  #10 
a = 8'd99; b = 8'd142;  #10 
a = 8'd99; b = 8'd143;  #10 
a = 8'd99; b = 8'd144;  #10 
a = 8'd99; b = 8'd145;  #10 
a = 8'd99; b = 8'd146;  #10 
a = 8'd99; b = 8'd147;  #10 
a = 8'd99; b = 8'd148;  #10 
a = 8'd99; b = 8'd149;  #10 
a = 8'd99; b = 8'd150;  #10 
a = 8'd99; b = 8'd151;  #10 
a = 8'd99; b = 8'd152;  #10 
a = 8'd99; b = 8'd153;  #10 
a = 8'd99; b = 8'd154;  #10 
a = 8'd99; b = 8'd155;  #10 
a = 8'd99; b = 8'd156;  #10 
a = 8'd99; b = 8'd157;  #10 
a = 8'd99; b = 8'd158;  #10 
a = 8'd99; b = 8'd159;  #10 
a = 8'd99; b = 8'd160;  #10 
a = 8'd99; b = 8'd161;  #10 
a = 8'd99; b = 8'd162;  #10 
a = 8'd99; b = 8'd163;  #10 
a = 8'd99; b = 8'd164;  #10 
a = 8'd99; b = 8'd165;  #10 
a = 8'd99; b = 8'd166;  #10 
a = 8'd99; b = 8'd167;  #10 
a = 8'd99; b = 8'd168;  #10 
a = 8'd99; b = 8'd169;  #10 
a = 8'd99; b = 8'd170;  #10 
a = 8'd99; b = 8'd171;  #10 
a = 8'd99; b = 8'd172;  #10 
a = 8'd99; b = 8'd173;  #10 
a = 8'd99; b = 8'd174;  #10 
a = 8'd99; b = 8'd175;  #10 
a = 8'd99; b = 8'd176;  #10 
a = 8'd99; b = 8'd177;  #10 
a = 8'd99; b = 8'd178;  #10 
a = 8'd99; b = 8'd179;  #10 
a = 8'd99; b = 8'd180;  #10 
a = 8'd99; b = 8'd181;  #10 
a = 8'd99; b = 8'd182;  #10 
a = 8'd99; b = 8'd183;  #10 
a = 8'd99; b = 8'd184;  #10 
a = 8'd99; b = 8'd185;  #10 
a = 8'd99; b = 8'd186;  #10 
a = 8'd99; b = 8'd187;  #10 
a = 8'd99; b = 8'd188;  #10 
a = 8'd99; b = 8'd189;  #10 
a = 8'd99; b = 8'd190;  #10 
a = 8'd99; b = 8'd191;  #10 
a = 8'd99; b = 8'd192;  #10 
a = 8'd99; b = 8'd193;  #10 
a = 8'd99; b = 8'd194;  #10 
a = 8'd99; b = 8'd195;  #10 
a = 8'd99; b = 8'd196;  #10 
a = 8'd99; b = 8'd197;  #10 
a = 8'd99; b = 8'd198;  #10 
a = 8'd99; b = 8'd199;  #10 
a = 8'd99; b = 8'd200;  #10 
a = 8'd99; b = 8'd201;  #10 
a = 8'd99; b = 8'd202;  #10 
a = 8'd99; b = 8'd203;  #10 
a = 8'd99; b = 8'd204;  #10 
a = 8'd99; b = 8'd205;  #10 
a = 8'd99; b = 8'd206;  #10 
a = 8'd99; b = 8'd207;  #10 
a = 8'd99; b = 8'd208;  #10 
a = 8'd99; b = 8'd209;  #10 
a = 8'd99; b = 8'd210;  #10 
a = 8'd99; b = 8'd211;  #10 
a = 8'd99; b = 8'd212;  #10 
a = 8'd99; b = 8'd213;  #10 
a = 8'd99; b = 8'd214;  #10 
a = 8'd99; b = 8'd215;  #10 
a = 8'd99; b = 8'd216;  #10 
a = 8'd99; b = 8'd217;  #10 
a = 8'd99; b = 8'd218;  #10 
a = 8'd99; b = 8'd219;  #10 
a = 8'd99; b = 8'd220;  #10 
a = 8'd99; b = 8'd221;  #10 
a = 8'd99; b = 8'd222;  #10 
a = 8'd99; b = 8'd223;  #10 
a = 8'd99; b = 8'd224;  #10 
a = 8'd99; b = 8'd225;  #10 
a = 8'd99; b = 8'd226;  #10 
a = 8'd99; b = 8'd227;  #10 
a = 8'd99; b = 8'd228;  #10 
a = 8'd99; b = 8'd229;  #10 
a = 8'd99; b = 8'd230;  #10 
a = 8'd99; b = 8'd231;  #10 
a = 8'd99; b = 8'd232;  #10 
a = 8'd99; b = 8'd233;  #10 
a = 8'd99; b = 8'd234;  #10 
a = 8'd99; b = 8'd235;  #10 
a = 8'd99; b = 8'd236;  #10 
a = 8'd99; b = 8'd237;  #10 
a = 8'd99; b = 8'd238;  #10 
a = 8'd99; b = 8'd239;  #10 
a = 8'd99; b = 8'd240;  #10 
a = 8'd99; b = 8'd241;  #10 
a = 8'd99; b = 8'd242;  #10 
a = 8'd99; b = 8'd243;  #10 
a = 8'd99; b = 8'd244;  #10 
a = 8'd99; b = 8'd245;  #10 
a = 8'd99; b = 8'd246;  #10 
a = 8'd99; b = 8'd247;  #10 
a = 8'd99; b = 8'd248;  #10 
a = 8'd99; b = 8'd249;  #10 
a = 8'd99; b = 8'd250;  #10 
a = 8'd99; b = 8'd251;  #10 
a = 8'd99; b = 8'd252;  #10 
a = 8'd99; b = 8'd253;  #10 
a = 8'd99; b = 8'd254;  #10 
a = 8'd99; b = 8'd255;  #10 
a = 8'd100; b = 8'd0;  #10 
a = 8'd100; b = 8'd1;  #10 
a = 8'd100; b = 8'd2;  #10 
a = 8'd100; b = 8'd3;  #10 
a = 8'd100; b = 8'd4;  #10 
a = 8'd100; b = 8'd5;  #10 
a = 8'd100; b = 8'd6;  #10 
a = 8'd100; b = 8'd7;  #10 
a = 8'd100; b = 8'd8;  #10 
a = 8'd100; b = 8'd9;  #10 
a = 8'd100; b = 8'd10;  #10 
a = 8'd100; b = 8'd11;  #10 
a = 8'd100; b = 8'd12;  #10 
a = 8'd100; b = 8'd13;  #10 
a = 8'd100; b = 8'd14;  #10 
a = 8'd100; b = 8'd15;  #10 
a = 8'd100; b = 8'd16;  #10 
a = 8'd100; b = 8'd17;  #10 
a = 8'd100; b = 8'd18;  #10 
a = 8'd100; b = 8'd19;  #10 
a = 8'd100; b = 8'd20;  #10 
a = 8'd100; b = 8'd21;  #10 
a = 8'd100; b = 8'd22;  #10 
a = 8'd100; b = 8'd23;  #10 
a = 8'd100; b = 8'd24;  #10 
a = 8'd100; b = 8'd25;  #10 
a = 8'd100; b = 8'd26;  #10 
a = 8'd100; b = 8'd27;  #10 
a = 8'd100; b = 8'd28;  #10 
a = 8'd100; b = 8'd29;  #10 
a = 8'd100; b = 8'd30;  #10 
a = 8'd100; b = 8'd31;  #10 
a = 8'd100; b = 8'd32;  #10 
a = 8'd100; b = 8'd33;  #10 
a = 8'd100; b = 8'd34;  #10 
a = 8'd100; b = 8'd35;  #10 
a = 8'd100; b = 8'd36;  #10 
a = 8'd100; b = 8'd37;  #10 
a = 8'd100; b = 8'd38;  #10 
a = 8'd100; b = 8'd39;  #10 
a = 8'd100; b = 8'd40;  #10 
a = 8'd100; b = 8'd41;  #10 
a = 8'd100; b = 8'd42;  #10 
a = 8'd100; b = 8'd43;  #10 
a = 8'd100; b = 8'd44;  #10 
a = 8'd100; b = 8'd45;  #10 
a = 8'd100; b = 8'd46;  #10 
a = 8'd100; b = 8'd47;  #10 
a = 8'd100; b = 8'd48;  #10 
a = 8'd100; b = 8'd49;  #10 
a = 8'd100; b = 8'd50;  #10 
a = 8'd100; b = 8'd51;  #10 
a = 8'd100; b = 8'd52;  #10 
a = 8'd100; b = 8'd53;  #10 
a = 8'd100; b = 8'd54;  #10 
a = 8'd100; b = 8'd55;  #10 
a = 8'd100; b = 8'd56;  #10 
a = 8'd100; b = 8'd57;  #10 
a = 8'd100; b = 8'd58;  #10 
a = 8'd100; b = 8'd59;  #10 
a = 8'd100; b = 8'd60;  #10 
a = 8'd100; b = 8'd61;  #10 
a = 8'd100; b = 8'd62;  #10 
a = 8'd100; b = 8'd63;  #10 
a = 8'd100; b = 8'd64;  #10 
a = 8'd100; b = 8'd65;  #10 
a = 8'd100; b = 8'd66;  #10 
a = 8'd100; b = 8'd67;  #10 
a = 8'd100; b = 8'd68;  #10 
a = 8'd100; b = 8'd69;  #10 
a = 8'd100; b = 8'd70;  #10 
a = 8'd100; b = 8'd71;  #10 
a = 8'd100; b = 8'd72;  #10 
a = 8'd100; b = 8'd73;  #10 
a = 8'd100; b = 8'd74;  #10 
a = 8'd100; b = 8'd75;  #10 
a = 8'd100; b = 8'd76;  #10 
a = 8'd100; b = 8'd77;  #10 
a = 8'd100; b = 8'd78;  #10 
a = 8'd100; b = 8'd79;  #10 
a = 8'd100; b = 8'd80;  #10 
a = 8'd100; b = 8'd81;  #10 
a = 8'd100; b = 8'd82;  #10 
a = 8'd100; b = 8'd83;  #10 
a = 8'd100; b = 8'd84;  #10 
a = 8'd100; b = 8'd85;  #10 
a = 8'd100; b = 8'd86;  #10 
a = 8'd100; b = 8'd87;  #10 
a = 8'd100; b = 8'd88;  #10 
a = 8'd100; b = 8'd89;  #10 
a = 8'd100; b = 8'd90;  #10 
a = 8'd100; b = 8'd91;  #10 
a = 8'd100; b = 8'd92;  #10 
a = 8'd100; b = 8'd93;  #10 
a = 8'd100; b = 8'd94;  #10 
a = 8'd100; b = 8'd95;  #10 
a = 8'd100; b = 8'd96;  #10 
a = 8'd100; b = 8'd97;  #10 
a = 8'd100; b = 8'd98;  #10 
a = 8'd100; b = 8'd99;  #10 
a = 8'd100; b = 8'd100;  #10 
a = 8'd100; b = 8'd101;  #10 
a = 8'd100; b = 8'd102;  #10 
a = 8'd100; b = 8'd103;  #10 
a = 8'd100; b = 8'd104;  #10 
a = 8'd100; b = 8'd105;  #10 
a = 8'd100; b = 8'd106;  #10 
a = 8'd100; b = 8'd107;  #10 
a = 8'd100; b = 8'd108;  #10 
a = 8'd100; b = 8'd109;  #10 
a = 8'd100; b = 8'd110;  #10 
a = 8'd100; b = 8'd111;  #10 
a = 8'd100; b = 8'd112;  #10 
a = 8'd100; b = 8'd113;  #10 
a = 8'd100; b = 8'd114;  #10 
a = 8'd100; b = 8'd115;  #10 
a = 8'd100; b = 8'd116;  #10 
a = 8'd100; b = 8'd117;  #10 
a = 8'd100; b = 8'd118;  #10 
a = 8'd100; b = 8'd119;  #10 
a = 8'd100; b = 8'd120;  #10 
a = 8'd100; b = 8'd121;  #10 
a = 8'd100; b = 8'd122;  #10 
a = 8'd100; b = 8'd123;  #10 
a = 8'd100; b = 8'd124;  #10 
a = 8'd100; b = 8'd125;  #10 
a = 8'd100; b = 8'd126;  #10 
a = 8'd100; b = 8'd127;  #10 
a = 8'd100; b = 8'd128;  #10 
a = 8'd100; b = 8'd129;  #10 
a = 8'd100; b = 8'd130;  #10 
a = 8'd100; b = 8'd131;  #10 
a = 8'd100; b = 8'd132;  #10 
a = 8'd100; b = 8'd133;  #10 
a = 8'd100; b = 8'd134;  #10 
a = 8'd100; b = 8'd135;  #10 
a = 8'd100; b = 8'd136;  #10 
a = 8'd100; b = 8'd137;  #10 
a = 8'd100; b = 8'd138;  #10 
a = 8'd100; b = 8'd139;  #10 
a = 8'd100; b = 8'd140;  #10 
a = 8'd100; b = 8'd141;  #10 
a = 8'd100; b = 8'd142;  #10 
a = 8'd100; b = 8'd143;  #10 
a = 8'd100; b = 8'd144;  #10 
a = 8'd100; b = 8'd145;  #10 
a = 8'd100; b = 8'd146;  #10 
a = 8'd100; b = 8'd147;  #10 
a = 8'd100; b = 8'd148;  #10 
a = 8'd100; b = 8'd149;  #10 
a = 8'd100; b = 8'd150;  #10 
a = 8'd100; b = 8'd151;  #10 
a = 8'd100; b = 8'd152;  #10 
a = 8'd100; b = 8'd153;  #10 
a = 8'd100; b = 8'd154;  #10 
a = 8'd100; b = 8'd155;  #10 
a = 8'd100; b = 8'd156;  #10 
a = 8'd100; b = 8'd157;  #10 
a = 8'd100; b = 8'd158;  #10 
a = 8'd100; b = 8'd159;  #10 
a = 8'd100; b = 8'd160;  #10 
a = 8'd100; b = 8'd161;  #10 
a = 8'd100; b = 8'd162;  #10 
a = 8'd100; b = 8'd163;  #10 
a = 8'd100; b = 8'd164;  #10 
a = 8'd100; b = 8'd165;  #10 
a = 8'd100; b = 8'd166;  #10 
a = 8'd100; b = 8'd167;  #10 
a = 8'd100; b = 8'd168;  #10 
a = 8'd100; b = 8'd169;  #10 
a = 8'd100; b = 8'd170;  #10 
a = 8'd100; b = 8'd171;  #10 
a = 8'd100; b = 8'd172;  #10 
a = 8'd100; b = 8'd173;  #10 
a = 8'd100; b = 8'd174;  #10 
a = 8'd100; b = 8'd175;  #10 
a = 8'd100; b = 8'd176;  #10 
a = 8'd100; b = 8'd177;  #10 
a = 8'd100; b = 8'd178;  #10 
a = 8'd100; b = 8'd179;  #10 
a = 8'd100; b = 8'd180;  #10 
a = 8'd100; b = 8'd181;  #10 
a = 8'd100; b = 8'd182;  #10 
a = 8'd100; b = 8'd183;  #10 
a = 8'd100; b = 8'd184;  #10 
a = 8'd100; b = 8'd185;  #10 
a = 8'd100; b = 8'd186;  #10 
a = 8'd100; b = 8'd187;  #10 
a = 8'd100; b = 8'd188;  #10 
a = 8'd100; b = 8'd189;  #10 
a = 8'd100; b = 8'd190;  #10 
a = 8'd100; b = 8'd191;  #10 
a = 8'd100; b = 8'd192;  #10 
a = 8'd100; b = 8'd193;  #10 
a = 8'd100; b = 8'd194;  #10 
a = 8'd100; b = 8'd195;  #10 
a = 8'd100; b = 8'd196;  #10 
a = 8'd100; b = 8'd197;  #10 
a = 8'd100; b = 8'd198;  #10 
a = 8'd100; b = 8'd199;  #10 
a = 8'd100; b = 8'd200;  #10 
a = 8'd100; b = 8'd201;  #10 
a = 8'd100; b = 8'd202;  #10 
a = 8'd100; b = 8'd203;  #10 
a = 8'd100; b = 8'd204;  #10 
a = 8'd100; b = 8'd205;  #10 
a = 8'd100; b = 8'd206;  #10 
a = 8'd100; b = 8'd207;  #10 
a = 8'd100; b = 8'd208;  #10 
a = 8'd100; b = 8'd209;  #10 
a = 8'd100; b = 8'd210;  #10 
a = 8'd100; b = 8'd211;  #10 
a = 8'd100; b = 8'd212;  #10 
a = 8'd100; b = 8'd213;  #10 
a = 8'd100; b = 8'd214;  #10 
a = 8'd100; b = 8'd215;  #10 
a = 8'd100; b = 8'd216;  #10 
a = 8'd100; b = 8'd217;  #10 
a = 8'd100; b = 8'd218;  #10 
a = 8'd100; b = 8'd219;  #10 
a = 8'd100; b = 8'd220;  #10 
a = 8'd100; b = 8'd221;  #10 
a = 8'd100; b = 8'd222;  #10 
a = 8'd100; b = 8'd223;  #10 
a = 8'd100; b = 8'd224;  #10 
a = 8'd100; b = 8'd225;  #10 
a = 8'd100; b = 8'd226;  #10 
a = 8'd100; b = 8'd227;  #10 
a = 8'd100; b = 8'd228;  #10 
a = 8'd100; b = 8'd229;  #10 
a = 8'd100; b = 8'd230;  #10 
a = 8'd100; b = 8'd231;  #10 
a = 8'd100; b = 8'd232;  #10 
a = 8'd100; b = 8'd233;  #10 
a = 8'd100; b = 8'd234;  #10 
a = 8'd100; b = 8'd235;  #10 
a = 8'd100; b = 8'd236;  #10 
a = 8'd100; b = 8'd237;  #10 
a = 8'd100; b = 8'd238;  #10 
a = 8'd100; b = 8'd239;  #10 
a = 8'd100; b = 8'd240;  #10 
a = 8'd100; b = 8'd241;  #10 
a = 8'd100; b = 8'd242;  #10 
a = 8'd100; b = 8'd243;  #10 
a = 8'd100; b = 8'd244;  #10 
a = 8'd100; b = 8'd245;  #10 
a = 8'd100; b = 8'd246;  #10 
a = 8'd100; b = 8'd247;  #10 
a = 8'd100; b = 8'd248;  #10 
a = 8'd100; b = 8'd249;  #10 
a = 8'd100; b = 8'd250;  #10 
a = 8'd100; b = 8'd251;  #10 
a = 8'd100; b = 8'd252;  #10 
a = 8'd100; b = 8'd253;  #10 
a = 8'd100; b = 8'd254;  #10 
a = 8'd100; b = 8'd255;  #10 
a = 8'd101; b = 8'd0;  #10 
a = 8'd101; b = 8'd1;  #10 
a = 8'd101; b = 8'd2;  #10 
a = 8'd101; b = 8'd3;  #10 
a = 8'd101; b = 8'd4;  #10 
a = 8'd101; b = 8'd5;  #10 
a = 8'd101; b = 8'd6;  #10 
a = 8'd101; b = 8'd7;  #10 
a = 8'd101; b = 8'd8;  #10 
a = 8'd101; b = 8'd9;  #10 
a = 8'd101; b = 8'd10;  #10 
a = 8'd101; b = 8'd11;  #10 
a = 8'd101; b = 8'd12;  #10 
a = 8'd101; b = 8'd13;  #10 
a = 8'd101; b = 8'd14;  #10 
a = 8'd101; b = 8'd15;  #10 
a = 8'd101; b = 8'd16;  #10 
a = 8'd101; b = 8'd17;  #10 
a = 8'd101; b = 8'd18;  #10 
a = 8'd101; b = 8'd19;  #10 
a = 8'd101; b = 8'd20;  #10 
a = 8'd101; b = 8'd21;  #10 
a = 8'd101; b = 8'd22;  #10 
a = 8'd101; b = 8'd23;  #10 
a = 8'd101; b = 8'd24;  #10 
a = 8'd101; b = 8'd25;  #10 
a = 8'd101; b = 8'd26;  #10 
a = 8'd101; b = 8'd27;  #10 
a = 8'd101; b = 8'd28;  #10 
a = 8'd101; b = 8'd29;  #10 
a = 8'd101; b = 8'd30;  #10 
a = 8'd101; b = 8'd31;  #10 
a = 8'd101; b = 8'd32;  #10 
a = 8'd101; b = 8'd33;  #10 
a = 8'd101; b = 8'd34;  #10 
a = 8'd101; b = 8'd35;  #10 
a = 8'd101; b = 8'd36;  #10 
a = 8'd101; b = 8'd37;  #10 
a = 8'd101; b = 8'd38;  #10 
a = 8'd101; b = 8'd39;  #10 
a = 8'd101; b = 8'd40;  #10 
a = 8'd101; b = 8'd41;  #10 
a = 8'd101; b = 8'd42;  #10 
a = 8'd101; b = 8'd43;  #10 
a = 8'd101; b = 8'd44;  #10 
a = 8'd101; b = 8'd45;  #10 
a = 8'd101; b = 8'd46;  #10 
a = 8'd101; b = 8'd47;  #10 
a = 8'd101; b = 8'd48;  #10 
a = 8'd101; b = 8'd49;  #10 
a = 8'd101; b = 8'd50;  #10 
a = 8'd101; b = 8'd51;  #10 
a = 8'd101; b = 8'd52;  #10 
a = 8'd101; b = 8'd53;  #10 
a = 8'd101; b = 8'd54;  #10 
a = 8'd101; b = 8'd55;  #10 
a = 8'd101; b = 8'd56;  #10 
a = 8'd101; b = 8'd57;  #10 
a = 8'd101; b = 8'd58;  #10 
a = 8'd101; b = 8'd59;  #10 
a = 8'd101; b = 8'd60;  #10 
a = 8'd101; b = 8'd61;  #10 
a = 8'd101; b = 8'd62;  #10 
a = 8'd101; b = 8'd63;  #10 
a = 8'd101; b = 8'd64;  #10 
a = 8'd101; b = 8'd65;  #10 
a = 8'd101; b = 8'd66;  #10 
a = 8'd101; b = 8'd67;  #10 
a = 8'd101; b = 8'd68;  #10 
a = 8'd101; b = 8'd69;  #10 
a = 8'd101; b = 8'd70;  #10 
a = 8'd101; b = 8'd71;  #10 
a = 8'd101; b = 8'd72;  #10 
a = 8'd101; b = 8'd73;  #10 
a = 8'd101; b = 8'd74;  #10 
a = 8'd101; b = 8'd75;  #10 
a = 8'd101; b = 8'd76;  #10 
a = 8'd101; b = 8'd77;  #10 
a = 8'd101; b = 8'd78;  #10 
a = 8'd101; b = 8'd79;  #10 
a = 8'd101; b = 8'd80;  #10 
a = 8'd101; b = 8'd81;  #10 
a = 8'd101; b = 8'd82;  #10 
a = 8'd101; b = 8'd83;  #10 
a = 8'd101; b = 8'd84;  #10 
a = 8'd101; b = 8'd85;  #10 
a = 8'd101; b = 8'd86;  #10 
a = 8'd101; b = 8'd87;  #10 
a = 8'd101; b = 8'd88;  #10 
a = 8'd101; b = 8'd89;  #10 
a = 8'd101; b = 8'd90;  #10 
a = 8'd101; b = 8'd91;  #10 
a = 8'd101; b = 8'd92;  #10 
a = 8'd101; b = 8'd93;  #10 
a = 8'd101; b = 8'd94;  #10 
a = 8'd101; b = 8'd95;  #10 
a = 8'd101; b = 8'd96;  #10 
a = 8'd101; b = 8'd97;  #10 
a = 8'd101; b = 8'd98;  #10 
a = 8'd101; b = 8'd99;  #10 
a = 8'd101; b = 8'd100;  #10 
a = 8'd101; b = 8'd101;  #10 
a = 8'd101; b = 8'd102;  #10 
a = 8'd101; b = 8'd103;  #10 
a = 8'd101; b = 8'd104;  #10 
a = 8'd101; b = 8'd105;  #10 
a = 8'd101; b = 8'd106;  #10 
a = 8'd101; b = 8'd107;  #10 
a = 8'd101; b = 8'd108;  #10 
a = 8'd101; b = 8'd109;  #10 
a = 8'd101; b = 8'd110;  #10 
a = 8'd101; b = 8'd111;  #10 
a = 8'd101; b = 8'd112;  #10 
a = 8'd101; b = 8'd113;  #10 
a = 8'd101; b = 8'd114;  #10 
a = 8'd101; b = 8'd115;  #10 
a = 8'd101; b = 8'd116;  #10 
a = 8'd101; b = 8'd117;  #10 
a = 8'd101; b = 8'd118;  #10 
a = 8'd101; b = 8'd119;  #10 
a = 8'd101; b = 8'd120;  #10 
a = 8'd101; b = 8'd121;  #10 
a = 8'd101; b = 8'd122;  #10 
a = 8'd101; b = 8'd123;  #10 
a = 8'd101; b = 8'd124;  #10 
a = 8'd101; b = 8'd125;  #10 
a = 8'd101; b = 8'd126;  #10 
a = 8'd101; b = 8'd127;  #10 
a = 8'd101; b = 8'd128;  #10 
a = 8'd101; b = 8'd129;  #10 
a = 8'd101; b = 8'd130;  #10 
a = 8'd101; b = 8'd131;  #10 
a = 8'd101; b = 8'd132;  #10 
a = 8'd101; b = 8'd133;  #10 
a = 8'd101; b = 8'd134;  #10 
a = 8'd101; b = 8'd135;  #10 
a = 8'd101; b = 8'd136;  #10 
a = 8'd101; b = 8'd137;  #10 
a = 8'd101; b = 8'd138;  #10 
a = 8'd101; b = 8'd139;  #10 
a = 8'd101; b = 8'd140;  #10 
a = 8'd101; b = 8'd141;  #10 
a = 8'd101; b = 8'd142;  #10 
a = 8'd101; b = 8'd143;  #10 
a = 8'd101; b = 8'd144;  #10 
a = 8'd101; b = 8'd145;  #10 
a = 8'd101; b = 8'd146;  #10 
a = 8'd101; b = 8'd147;  #10 
a = 8'd101; b = 8'd148;  #10 
a = 8'd101; b = 8'd149;  #10 
a = 8'd101; b = 8'd150;  #10 
a = 8'd101; b = 8'd151;  #10 
a = 8'd101; b = 8'd152;  #10 
a = 8'd101; b = 8'd153;  #10 
a = 8'd101; b = 8'd154;  #10 
a = 8'd101; b = 8'd155;  #10 
a = 8'd101; b = 8'd156;  #10 
a = 8'd101; b = 8'd157;  #10 
a = 8'd101; b = 8'd158;  #10 
a = 8'd101; b = 8'd159;  #10 
a = 8'd101; b = 8'd160;  #10 
a = 8'd101; b = 8'd161;  #10 
a = 8'd101; b = 8'd162;  #10 
a = 8'd101; b = 8'd163;  #10 
a = 8'd101; b = 8'd164;  #10 
a = 8'd101; b = 8'd165;  #10 
a = 8'd101; b = 8'd166;  #10 
a = 8'd101; b = 8'd167;  #10 
a = 8'd101; b = 8'd168;  #10 
a = 8'd101; b = 8'd169;  #10 
a = 8'd101; b = 8'd170;  #10 
a = 8'd101; b = 8'd171;  #10 
a = 8'd101; b = 8'd172;  #10 
a = 8'd101; b = 8'd173;  #10 
a = 8'd101; b = 8'd174;  #10 
a = 8'd101; b = 8'd175;  #10 
a = 8'd101; b = 8'd176;  #10 
a = 8'd101; b = 8'd177;  #10 
a = 8'd101; b = 8'd178;  #10 
a = 8'd101; b = 8'd179;  #10 
a = 8'd101; b = 8'd180;  #10 
a = 8'd101; b = 8'd181;  #10 
a = 8'd101; b = 8'd182;  #10 
a = 8'd101; b = 8'd183;  #10 
a = 8'd101; b = 8'd184;  #10 
a = 8'd101; b = 8'd185;  #10 
a = 8'd101; b = 8'd186;  #10 
a = 8'd101; b = 8'd187;  #10 
a = 8'd101; b = 8'd188;  #10 
a = 8'd101; b = 8'd189;  #10 
a = 8'd101; b = 8'd190;  #10 
a = 8'd101; b = 8'd191;  #10 
a = 8'd101; b = 8'd192;  #10 
a = 8'd101; b = 8'd193;  #10 
a = 8'd101; b = 8'd194;  #10 
a = 8'd101; b = 8'd195;  #10 
a = 8'd101; b = 8'd196;  #10 
a = 8'd101; b = 8'd197;  #10 
a = 8'd101; b = 8'd198;  #10 
a = 8'd101; b = 8'd199;  #10 
a = 8'd101; b = 8'd200;  #10 
a = 8'd101; b = 8'd201;  #10 
a = 8'd101; b = 8'd202;  #10 
a = 8'd101; b = 8'd203;  #10 
a = 8'd101; b = 8'd204;  #10 
a = 8'd101; b = 8'd205;  #10 
a = 8'd101; b = 8'd206;  #10 
a = 8'd101; b = 8'd207;  #10 
a = 8'd101; b = 8'd208;  #10 
a = 8'd101; b = 8'd209;  #10 
a = 8'd101; b = 8'd210;  #10 
a = 8'd101; b = 8'd211;  #10 
a = 8'd101; b = 8'd212;  #10 
a = 8'd101; b = 8'd213;  #10 
a = 8'd101; b = 8'd214;  #10 
a = 8'd101; b = 8'd215;  #10 
a = 8'd101; b = 8'd216;  #10 
a = 8'd101; b = 8'd217;  #10 
a = 8'd101; b = 8'd218;  #10 
a = 8'd101; b = 8'd219;  #10 
a = 8'd101; b = 8'd220;  #10 
a = 8'd101; b = 8'd221;  #10 
a = 8'd101; b = 8'd222;  #10 
a = 8'd101; b = 8'd223;  #10 
a = 8'd101; b = 8'd224;  #10 
a = 8'd101; b = 8'd225;  #10 
a = 8'd101; b = 8'd226;  #10 
a = 8'd101; b = 8'd227;  #10 
a = 8'd101; b = 8'd228;  #10 
a = 8'd101; b = 8'd229;  #10 
a = 8'd101; b = 8'd230;  #10 
a = 8'd101; b = 8'd231;  #10 
a = 8'd101; b = 8'd232;  #10 
a = 8'd101; b = 8'd233;  #10 
a = 8'd101; b = 8'd234;  #10 
a = 8'd101; b = 8'd235;  #10 
a = 8'd101; b = 8'd236;  #10 
a = 8'd101; b = 8'd237;  #10 
a = 8'd101; b = 8'd238;  #10 
a = 8'd101; b = 8'd239;  #10 
a = 8'd101; b = 8'd240;  #10 
a = 8'd101; b = 8'd241;  #10 
a = 8'd101; b = 8'd242;  #10 
a = 8'd101; b = 8'd243;  #10 
a = 8'd101; b = 8'd244;  #10 
a = 8'd101; b = 8'd245;  #10 
a = 8'd101; b = 8'd246;  #10 
a = 8'd101; b = 8'd247;  #10 
a = 8'd101; b = 8'd248;  #10 
a = 8'd101; b = 8'd249;  #10 
a = 8'd101; b = 8'd250;  #10 
a = 8'd101; b = 8'd251;  #10 
a = 8'd101; b = 8'd252;  #10 
a = 8'd101; b = 8'd253;  #10 
a = 8'd101; b = 8'd254;  #10 
a = 8'd101; b = 8'd255;  #10 
a = 8'd102; b = 8'd0;  #10 
a = 8'd102; b = 8'd1;  #10 
a = 8'd102; b = 8'd2;  #10 
a = 8'd102; b = 8'd3;  #10 
a = 8'd102; b = 8'd4;  #10 
a = 8'd102; b = 8'd5;  #10 
a = 8'd102; b = 8'd6;  #10 
a = 8'd102; b = 8'd7;  #10 
a = 8'd102; b = 8'd8;  #10 
a = 8'd102; b = 8'd9;  #10 
a = 8'd102; b = 8'd10;  #10 
a = 8'd102; b = 8'd11;  #10 
a = 8'd102; b = 8'd12;  #10 
a = 8'd102; b = 8'd13;  #10 
a = 8'd102; b = 8'd14;  #10 
a = 8'd102; b = 8'd15;  #10 
a = 8'd102; b = 8'd16;  #10 
a = 8'd102; b = 8'd17;  #10 
a = 8'd102; b = 8'd18;  #10 
a = 8'd102; b = 8'd19;  #10 
a = 8'd102; b = 8'd20;  #10 
a = 8'd102; b = 8'd21;  #10 
a = 8'd102; b = 8'd22;  #10 
a = 8'd102; b = 8'd23;  #10 
a = 8'd102; b = 8'd24;  #10 
a = 8'd102; b = 8'd25;  #10 
a = 8'd102; b = 8'd26;  #10 
a = 8'd102; b = 8'd27;  #10 
a = 8'd102; b = 8'd28;  #10 
a = 8'd102; b = 8'd29;  #10 
a = 8'd102; b = 8'd30;  #10 
a = 8'd102; b = 8'd31;  #10 
a = 8'd102; b = 8'd32;  #10 
a = 8'd102; b = 8'd33;  #10 
a = 8'd102; b = 8'd34;  #10 
a = 8'd102; b = 8'd35;  #10 
a = 8'd102; b = 8'd36;  #10 
a = 8'd102; b = 8'd37;  #10 
a = 8'd102; b = 8'd38;  #10 
a = 8'd102; b = 8'd39;  #10 
a = 8'd102; b = 8'd40;  #10 
a = 8'd102; b = 8'd41;  #10 
a = 8'd102; b = 8'd42;  #10 
a = 8'd102; b = 8'd43;  #10 
a = 8'd102; b = 8'd44;  #10 
a = 8'd102; b = 8'd45;  #10 
a = 8'd102; b = 8'd46;  #10 
a = 8'd102; b = 8'd47;  #10 
a = 8'd102; b = 8'd48;  #10 
a = 8'd102; b = 8'd49;  #10 
a = 8'd102; b = 8'd50;  #10 
a = 8'd102; b = 8'd51;  #10 
a = 8'd102; b = 8'd52;  #10 
a = 8'd102; b = 8'd53;  #10 
a = 8'd102; b = 8'd54;  #10 
a = 8'd102; b = 8'd55;  #10 
a = 8'd102; b = 8'd56;  #10 
a = 8'd102; b = 8'd57;  #10 
a = 8'd102; b = 8'd58;  #10 
a = 8'd102; b = 8'd59;  #10 
a = 8'd102; b = 8'd60;  #10 
a = 8'd102; b = 8'd61;  #10 
a = 8'd102; b = 8'd62;  #10 
a = 8'd102; b = 8'd63;  #10 
a = 8'd102; b = 8'd64;  #10 
a = 8'd102; b = 8'd65;  #10 
a = 8'd102; b = 8'd66;  #10 
a = 8'd102; b = 8'd67;  #10 
a = 8'd102; b = 8'd68;  #10 
a = 8'd102; b = 8'd69;  #10 
a = 8'd102; b = 8'd70;  #10 
a = 8'd102; b = 8'd71;  #10 
a = 8'd102; b = 8'd72;  #10 
a = 8'd102; b = 8'd73;  #10 
a = 8'd102; b = 8'd74;  #10 
a = 8'd102; b = 8'd75;  #10 
a = 8'd102; b = 8'd76;  #10 
a = 8'd102; b = 8'd77;  #10 
a = 8'd102; b = 8'd78;  #10 
a = 8'd102; b = 8'd79;  #10 
a = 8'd102; b = 8'd80;  #10 
a = 8'd102; b = 8'd81;  #10 
a = 8'd102; b = 8'd82;  #10 
a = 8'd102; b = 8'd83;  #10 
a = 8'd102; b = 8'd84;  #10 
a = 8'd102; b = 8'd85;  #10 
a = 8'd102; b = 8'd86;  #10 
a = 8'd102; b = 8'd87;  #10 
a = 8'd102; b = 8'd88;  #10 
a = 8'd102; b = 8'd89;  #10 
a = 8'd102; b = 8'd90;  #10 
a = 8'd102; b = 8'd91;  #10 
a = 8'd102; b = 8'd92;  #10 
a = 8'd102; b = 8'd93;  #10 
a = 8'd102; b = 8'd94;  #10 
a = 8'd102; b = 8'd95;  #10 
a = 8'd102; b = 8'd96;  #10 
a = 8'd102; b = 8'd97;  #10 
a = 8'd102; b = 8'd98;  #10 
a = 8'd102; b = 8'd99;  #10 
a = 8'd102; b = 8'd100;  #10 
a = 8'd102; b = 8'd101;  #10 
a = 8'd102; b = 8'd102;  #10 
a = 8'd102; b = 8'd103;  #10 
a = 8'd102; b = 8'd104;  #10 
a = 8'd102; b = 8'd105;  #10 
a = 8'd102; b = 8'd106;  #10 
a = 8'd102; b = 8'd107;  #10 
a = 8'd102; b = 8'd108;  #10 
a = 8'd102; b = 8'd109;  #10 
a = 8'd102; b = 8'd110;  #10 
a = 8'd102; b = 8'd111;  #10 
a = 8'd102; b = 8'd112;  #10 
a = 8'd102; b = 8'd113;  #10 
a = 8'd102; b = 8'd114;  #10 
a = 8'd102; b = 8'd115;  #10 
a = 8'd102; b = 8'd116;  #10 
a = 8'd102; b = 8'd117;  #10 
a = 8'd102; b = 8'd118;  #10 
a = 8'd102; b = 8'd119;  #10 
a = 8'd102; b = 8'd120;  #10 
a = 8'd102; b = 8'd121;  #10 
a = 8'd102; b = 8'd122;  #10 
a = 8'd102; b = 8'd123;  #10 
a = 8'd102; b = 8'd124;  #10 
a = 8'd102; b = 8'd125;  #10 
a = 8'd102; b = 8'd126;  #10 
a = 8'd102; b = 8'd127;  #10 
a = 8'd102; b = 8'd128;  #10 
a = 8'd102; b = 8'd129;  #10 
a = 8'd102; b = 8'd130;  #10 
a = 8'd102; b = 8'd131;  #10 
a = 8'd102; b = 8'd132;  #10 
a = 8'd102; b = 8'd133;  #10 
a = 8'd102; b = 8'd134;  #10 
a = 8'd102; b = 8'd135;  #10 
a = 8'd102; b = 8'd136;  #10 
a = 8'd102; b = 8'd137;  #10 
a = 8'd102; b = 8'd138;  #10 
a = 8'd102; b = 8'd139;  #10 
a = 8'd102; b = 8'd140;  #10 
a = 8'd102; b = 8'd141;  #10 
a = 8'd102; b = 8'd142;  #10 
a = 8'd102; b = 8'd143;  #10 
a = 8'd102; b = 8'd144;  #10 
a = 8'd102; b = 8'd145;  #10 
a = 8'd102; b = 8'd146;  #10 
a = 8'd102; b = 8'd147;  #10 
a = 8'd102; b = 8'd148;  #10 
a = 8'd102; b = 8'd149;  #10 
a = 8'd102; b = 8'd150;  #10 
a = 8'd102; b = 8'd151;  #10 
a = 8'd102; b = 8'd152;  #10 
a = 8'd102; b = 8'd153;  #10 
a = 8'd102; b = 8'd154;  #10 
a = 8'd102; b = 8'd155;  #10 
a = 8'd102; b = 8'd156;  #10 
a = 8'd102; b = 8'd157;  #10 
a = 8'd102; b = 8'd158;  #10 
a = 8'd102; b = 8'd159;  #10 
a = 8'd102; b = 8'd160;  #10 
a = 8'd102; b = 8'd161;  #10 
a = 8'd102; b = 8'd162;  #10 
a = 8'd102; b = 8'd163;  #10 
a = 8'd102; b = 8'd164;  #10 
a = 8'd102; b = 8'd165;  #10 
a = 8'd102; b = 8'd166;  #10 
a = 8'd102; b = 8'd167;  #10 
a = 8'd102; b = 8'd168;  #10 
a = 8'd102; b = 8'd169;  #10 
a = 8'd102; b = 8'd170;  #10 
a = 8'd102; b = 8'd171;  #10 
a = 8'd102; b = 8'd172;  #10 
a = 8'd102; b = 8'd173;  #10 
a = 8'd102; b = 8'd174;  #10 
a = 8'd102; b = 8'd175;  #10 
a = 8'd102; b = 8'd176;  #10 
a = 8'd102; b = 8'd177;  #10 
a = 8'd102; b = 8'd178;  #10 
a = 8'd102; b = 8'd179;  #10 
a = 8'd102; b = 8'd180;  #10 
a = 8'd102; b = 8'd181;  #10 
a = 8'd102; b = 8'd182;  #10 
a = 8'd102; b = 8'd183;  #10 
a = 8'd102; b = 8'd184;  #10 
a = 8'd102; b = 8'd185;  #10 
a = 8'd102; b = 8'd186;  #10 
a = 8'd102; b = 8'd187;  #10 
a = 8'd102; b = 8'd188;  #10 
a = 8'd102; b = 8'd189;  #10 
a = 8'd102; b = 8'd190;  #10 
a = 8'd102; b = 8'd191;  #10 
a = 8'd102; b = 8'd192;  #10 
a = 8'd102; b = 8'd193;  #10 
a = 8'd102; b = 8'd194;  #10 
a = 8'd102; b = 8'd195;  #10 
a = 8'd102; b = 8'd196;  #10 
a = 8'd102; b = 8'd197;  #10 
a = 8'd102; b = 8'd198;  #10 
a = 8'd102; b = 8'd199;  #10 
a = 8'd102; b = 8'd200;  #10 
a = 8'd102; b = 8'd201;  #10 
a = 8'd102; b = 8'd202;  #10 
a = 8'd102; b = 8'd203;  #10 
a = 8'd102; b = 8'd204;  #10 
a = 8'd102; b = 8'd205;  #10 
a = 8'd102; b = 8'd206;  #10 
a = 8'd102; b = 8'd207;  #10 
a = 8'd102; b = 8'd208;  #10 
a = 8'd102; b = 8'd209;  #10 
a = 8'd102; b = 8'd210;  #10 
a = 8'd102; b = 8'd211;  #10 
a = 8'd102; b = 8'd212;  #10 
a = 8'd102; b = 8'd213;  #10 
a = 8'd102; b = 8'd214;  #10 
a = 8'd102; b = 8'd215;  #10 
a = 8'd102; b = 8'd216;  #10 
a = 8'd102; b = 8'd217;  #10 
a = 8'd102; b = 8'd218;  #10 
a = 8'd102; b = 8'd219;  #10 
a = 8'd102; b = 8'd220;  #10 
a = 8'd102; b = 8'd221;  #10 
a = 8'd102; b = 8'd222;  #10 
a = 8'd102; b = 8'd223;  #10 
a = 8'd102; b = 8'd224;  #10 
a = 8'd102; b = 8'd225;  #10 
a = 8'd102; b = 8'd226;  #10 
a = 8'd102; b = 8'd227;  #10 
a = 8'd102; b = 8'd228;  #10 
a = 8'd102; b = 8'd229;  #10 
a = 8'd102; b = 8'd230;  #10 
a = 8'd102; b = 8'd231;  #10 
a = 8'd102; b = 8'd232;  #10 
a = 8'd102; b = 8'd233;  #10 
a = 8'd102; b = 8'd234;  #10 
a = 8'd102; b = 8'd235;  #10 
a = 8'd102; b = 8'd236;  #10 
a = 8'd102; b = 8'd237;  #10 
a = 8'd102; b = 8'd238;  #10 
a = 8'd102; b = 8'd239;  #10 
a = 8'd102; b = 8'd240;  #10 
a = 8'd102; b = 8'd241;  #10 
a = 8'd102; b = 8'd242;  #10 
a = 8'd102; b = 8'd243;  #10 
a = 8'd102; b = 8'd244;  #10 
a = 8'd102; b = 8'd245;  #10 
a = 8'd102; b = 8'd246;  #10 
a = 8'd102; b = 8'd247;  #10 
a = 8'd102; b = 8'd248;  #10 
a = 8'd102; b = 8'd249;  #10 
a = 8'd102; b = 8'd250;  #10 
a = 8'd102; b = 8'd251;  #10 
a = 8'd102; b = 8'd252;  #10 
a = 8'd102; b = 8'd253;  #10 
a = 8'd102; b = 8'd254;  #10 
a = 8'd102; b = 8'd255;  #10 
a = 8'd103; b = 8'd0;  #10 
a = 8'd103; b = 8'd1;  #10 
a = 8'd103; b = 8'd2;  #10 
a = 8'd103; b = 8'd3;  #10 
a = 8'd103; b = 8'd4;  #10 
a = 8'd103; b = 8'd5;  #10 
a = 8'd103; b = 8'd6;  #10 
a = 8'd103; b = 8'd7;  #10 
a = 8'd103; b = 8'd8;  #10 
a = 8'd103; b = 8'd9;  #10 
a = 8'd103; b = 8'd10;  #10 
a = 8'd103; b = 8'd11;  #10 
a = 8'd103; b = 8'd12;  #10 
a = 8'd103; b = 8'd13;  #10 
a = 8'd103; b = 8'd14;  #10 
a = 8'd103; b = 8'd15;  #10 
a = 8'd103; b = 8'd16;  #10 
a = 8'd103; b = 8'd17;  #10 
a = 8'd103; b = 8'd18;  #10 
a = 8'd103; b = 8'd19;  #10 
a = 8'd103; b = 8'd20;  #10 
a = 8'd103; b = 8'd21;  #10 
a = 8'd103; b = 8'd22;  #10 
a = 8'd103; b = 8'd23;  #10 
a = 8'd103; b = 8'd24;  #10 
a = 8'd103; b = 8'd25;  #10 
a = 8'd103; b = 8'd26;  #10 
a = 8'd103; b = 8'd27;  #10 
a = 8'd103; b = 8'd28;  #10 
a = 8'd103; b = 8'd29;  #10 
a = 8'd103; b = 8'd30;  #10 
a = 8'd103; b = 8'd31;  #10 
a = 8'd103; b = 8'd32;  #10 
a = 8'd103; b = 8'd33;  #10 
a = 8'd103; b = 8'd34;  #10 
a = 8'd103; b = 8'd35;  #10 
a = 8'd103; b = 8'd36;  #10 
a = 8'd103; b = 8'd37;  #10 
a = 8'd103; b = 8'd38;  #10 
a = 8'd103; b = 8'd39;  #10 
a = 8'd103; b = 8'd40;  #10 
a = 8'd103; b = 8'd41;  #10 
a = 8'd103; b = 8'd42;  #10 
a = 8'd103; b = 8'd43;  #10 
a = 8'd103; b = 8'd44;  #10 
a = 8'd103; b = 8'd45;  #10 
a = 8'd103; b = 8'd46;  #10 
a = 8'd103; b = 8'd47;  #10 
a = 8'd103; b = 8'd48;  #10 
a = 8'd103; b = 8'd49;  #10 
a = 8'd103; b = 8'd50;  #10 
a = 8'd103; b = 8'd51;  #10 
a = 8'd103; b = 8'd52;  #10 
a = 8'd103; b = 8'd53;  #10 
a = 8'd103; b = 8'd54;  #10 
a = 8'd103; b = 8'd55;  #10 
a = 8'd103; b = 8'd56;  #10 
a = 8'd103; b = 8'd57;  #10 
a = 8'd103; b = 8'd58;  #10 
a = 8'd103; b = 8'd59;  #10 
a = 8'd103; b = 8'd60;  #10 
a = 8'd103; b = 8'd61;  #10 
a = 8'd103; b = 8'd62;  #10 
a = 8'd103; b = 8'd63;  #10 
a = 8'd103; b = 8'd64;  #10 
a = 8'd103; b = 8'd65;  #10 
a = 8'd103; b = 8'd66;  #10 
a = 8'd103; b = 8'd67;  #10 
a = 8'd103; b = 8'd68;  #10 
a = 8'd103; b = 8'd69;  #10 
a = 8'd103; b = 8'd70;  #10 
a = 8'd103; b = 8'd71;  #10 
a = 8'd103; b = 8'd72;  #10 
a = 8'd103; b = 8'd73;  #10 
a = 8'd103; b = 8'd74;  #10 
a = 8'd103; b = 8'd75;  #10 
a = 8'd103; b = 8'd76;  #10 
a = 8'd103; b = 8'd77;  #10 
a = 8'd103; b = 8'd78;  #10 
a = 8'd103; b = 8'd79;  #10 
a = 8'd103; b = 8'd80;  #10 
a = 8'd103; b = 8'd81;  #10 
a = 8'd103; b = 8'd82;  #10 
a = 8'd103; b = 8'd83;  #10 
a = 8'd103; b = 8'd84;  #10 
a = 8'd103; b = 8'd85;  #10 
a = 8'd103; b = 8'd86;  #10 
a = 8'd103; b = 8'd87;  #10 
a = 8'd103; b = 8'd88;  #10 
a = 8'd103; b = 8'd89;  #10 
a = 8'd103; b = 8'd90;  #10 
a = 8'd103; b = 8'd91;  #10 
a = 8'd103; b = 8'd92;  #10 
a = 8'd103; b = 8'd93;  #10 
a = 8'd103; b = 8'd94;  #10 
a = 8'd103; b = 8'd95;  #10 
a = 8'd103; b = 8'd96;  #10 
a = 8'd103; b = 8'd97;  #10 
a = 8'd103; b = 8'd98;  #10 
a = 8'd103; b = 8'd99;  #10 
a = 8'd103; b = 8'd100;  #10 
a = 8'd103; b = 8'd101;  #10 
a = 8'd103; b = 8'd102;  #10 
a = 8'd103; b = 8'd103;  #10 
a = 8'd103; b = 8'd104;  #10 
a = 8'd103; b = 8'd105;  #10 
a = 8'd103; b = 8'd106;  #10 
a = 8'd103; b = 8'd107;  #10 
a = 8'd103; b = 8'd108;  #10 
a = 8'd103; b = 8'd109;  #10 
a = 8'd103; b = 8'd110;  #10 
a = 8'd103; b = 8'd111;  #10 
a = 8'd103; b = 8'd112;  #10 
a = 8'd103; b = 8'd113;  #10 
a = 8'd103; b = 8'd114;  #10 
a = 8'd103; b = 8'd115;  #10 
a = 8'd103; b = 8'd116;  #10 
a = 8'd103; b = 8'd117;  #10 
a = 8'd103; b = 8'd118;  #10 
a = 8'd103; b = 8'd119;  #10 
a = 8'd103; b = 8'd120;  #10 
a = 8'd103; b = 8'd121;  #10 
a = 8'd103; b = 8'd122;  #10 
a = 8'd103; b = 8'd123;  #10 
a = 8'd103; b = 8'd124;  #10 
a = 8'd103; b = 8'd125;  #10 
a = 8'd103; b = 8'd126;  #10 
a = 8'd103; b = 8'd127;  #10 
a = 8'd103; b = 8'd128;  #10 
a = 8'd103; b = 8'd129;  #10 
a = 8'd103; b = 8'd130;  #10 
a = 8'd103; b = 8'd131;  #10 
a = 8'd103; b = 8'd132;  #10 
a = 8'd103; b = 8'd133;  #10 
a = 8'd103; b = 8'd134;  #10 
a = 8'd103; b = 8'd135;  #10 
a = 8'd103; b = 8'd136;  #10 
a = 8'd103; b = 8'd137;  #10 
a = 8'd103; b = 8'd138;  #10 
a = 8'd103; b = 8'd139;  #10 
a = 8'd103; b = 8'd140;  #10 
a = 8'd103; b = 8'd141;  #10 
a = 8'd103; b = 8'd142;  #10 
a = 8'd103; b = 8'd143;  #10 
a = 8'd103; b = 8'd144;  #10 
a = 8'd103; b = 8'd145;  #10 
a = 8'd103; b = 8'd146;  #10 
a = 8'd103; b = 8'd147;  #10 
a = 8'd103; b = 8'd148;  #10 
a = 8'd103; b = 8'd149;  #10 
a = 8'd103; b = 8'd150;  #10 
a = 8'd103; b = 8'd151;  #10 
a = 8'd103; b = 8'd152;  #10 
a = 8'd103; b = 8'd153;  #10 
a = 8'd103; b = 8'd154;  #10 
a = 8'd103; b = 8'd155;  #10 
a = 8'd103; b = 8'd156;  #10 
a = 8'd103; b = 8'd157;  #10 
a = 8'd103; b = 8'd158;  #10 
a = 8'd103; b = 8'd159;  #10 
a = 8'd103; b = 8'd160;  #10 
a = 8'd103; b = 8'd161;  #10 
a = 8'd103; b = 8'd162;  #10 
a = 8'd103; b = 8'd163;  #10 
a = 8'd103; b = 8'd164;  #10 
a = 8'd103; b = 8'd165;  #10 
a = 8'd103; b = 8'd166;  #10 
a = 8'd103; b = 8'd167;  #10 
a = 8'd103; b = 8'd168;  #10 
a = 8'd103; b = 8'd169;  #10 
a = 8'd103; b = 8'd170;  #10 
a = 8'd103; b = 8'd171;  #10 
a = 8'd103; b = 8'd172;  #10 
a = 8'd103; b = 8'd173;  #10 
a = 8'd103; b = 8'd174;  #10 
a = 8'd103; b = 8'd175;  #10 
a = 8'd103; b = 8'd176;  #10 
a = 8'd103; b = 8'd177;  #10 
a = 8'd103; b = 8'd178;  #10 
a = 8'd103; b = 8'd179;  #10 
a = 8'd103; b = 8'd180;  #10 
a = 8'd103; b = 8'd181;  #10 
a = 8'd103; b = 8'd182;  #10 
a = 8'd103; b = 8'd183;  #10 
a = 8'd103; b = 8'd184;  #10 
a = 8'd103; b = 8'd185;  #10 
a = 8'd103; b = 8'd186;  #10 
a = 8'd103; b = 8'd187;  #10 
a = 8'd103; b = 8'd188;  #10 
a = 8'd103; b = 8'd189;  #10 
a = 8'd103; b = 8'd190;  #10 
a = 8'd103; b = 8'd191;  #10 
a = 8'd103; b = 8'd192;  #10 
a = 8'd103; b = 8'd193;  #10 
a = 8'd103; b = 8'd194;  #10 
a = 8'd103; b = 8'd195;  #10 
a = 8'd103; b = 8'd196;  #10 
a = 8'd103; b = 8'd197;  #10 
a = 8'd103; b = 8'd198;  #10 
a = 8'd103; b = 8'd199;  #10 
a = 8'd103; b = 8'd200;  #10 
a = 8'd103; b = 8'd201;  #10 
a = 8'd103; b = 8'd202;  #10 
a = 8'd103; b = 8'd203;  #10 
a = 8'd103; b = 8'd204;  #10 
a = 8'd103; b = 8'd205;  #10 
a = 8'd103; b = 8'd206;  #10 
a = 8'd103; b = 8'd207;  #10 
a = 8'd103; b = 8'd208;  #10 
a = 8'd103; b = 8'd209;  #10 
a = 8'd103; b = 8'd210;  #10 
a = 8'd103; b = 8'd211;  #10 
a = 8'd103; b = 8'd212;  #10 
a = 8'd103; b = 8'd213;  #10 
a = 8'd103; b = 8'd214;  #10 
a = 8'd103; b = 8'd215;  #10 
a = 8'd103; b = 8'd216;  #10 
a = 8'd103; b = 8'd217;  #10 
a = 8'd103; b = 8'd218;  #10 
a = 8'd103; b = 8'd219;  #10 
a = 8'd103; b = 8'd220;  #10 
a = 8'd103; b = 8'd221;  #10 
a = 8'd103; b = 8'd222;  #10 
a = 8'd103; b = 8'd223;  #10 
a = 8'd103; b = 8'd224;  #10 
a = 8'd103; b = 8'd225;  #10 
a = 8'd103; b = 8'd226;  #10 
a = 8'd103; b = 8'd227;  #10 
a = 8'd103; b = 8'd228;  #10 
a = 8'd103; b = 8'd229;  #10 
a = 8'd103; b = 8'd230;  #10 
a = 8'd103; b = 8'd231;  #10 
a = 8'd103; b = 8'd232;  #10 
a = 8'd103; b = 8'd233;  #10 
a = 8'd103; b = 8'd234;  #10 
a = 8'd103; b = 8'd235;  #10 
a = 8'd103; b = 8'd236;  #10 
a = 8'd103; b = 8'd237;  #10 
a = 8'd103; b = 8'd238;  #10 
a = 8'd103; b = 8'd239;  #10 
a = 8'd103; b = 8'd240;  #10 
a = 8'd103; b = 8'd241;  #10 
a = 8'd103; b = 8'd242;  #10 
a = 8'd103; b = 8'd243;  #10 
a = 8'd103; b = 8'd244;  #10 
a = 8'd103; b = 8'd245;  #10 
a = 8'd103; b = 8'd246;  #10 
a = 8'd103; b = 8'd247;  #10 
a = 8'd103; b = 8'd248;  #10 
a = 8'd103; b = 8'd249;  #10 
a = 8'd103; b = 8'd250;  #10 
a = 8'd103; b = 8'd251;  #10 
a = 8'd103; b = 8'd252;  #10 
a = 8'd103; b = 8'd253;  #10 
a = 8'd103; b = 8'd254;  #10 
a = 8'd103; b = 8'd255;  #10 
a = 8'd104; b = 8'd0;  #10 
a = 8'd104; b = 8'd1;  #10 
a = 8'd104; b = 8'd2;  #10 
a = 8'd104; b = 8'd3;  #10 
a = 8'd104; b = 8'd4;  #10 
a = 8'd104; b = 8'd5;  #10 
a = 8'd104; b = 8'd6;  #10 
a = 8'd104; b = 8'd7;  #10 
a = 8'd104; b = 8'd8;  #10 
a = 8'd104; b = 8'd9;  #10 
a = 8'd104; b = 8'd10;  #10 
a = 8'd104; b = 8'd11;  #10 
a = 8'd104; b = 8'd12;  #10 
a = 8'd104; b = 8'd13;  #10 
a = 8'd104; b = 8'd14;  #10 
a = 8'd104; b = 8'd15;  #10 
a = 8'd104; b = 8'd16;  #10 
a = 8'd104; b = 8'd17;  #10 
a = 8'd104; b = 8'd18;  #10 
a = 8'd104; b = 8'd19;  #10 
a = 8'd104; b = 8'd20;  #10 
a = 8'd104; b = 8'd21;  #10 
a = 8'd104; b = 8'd22;  #10 
a = 8'd104; b = 8'd23;  #10 
a = 8'd104; b = 8'd24;  #10 
a = 8'd104; b = 8'd25;  #10 
a = 8'd104; b = 8'd26;  #10 
a = 8'd104; b = 8'd27;  #10 
a = 8'd104; b = 8'd28;  #10 
a = 8'd104; b = 8'd29;  #10 
a = 8'd104; b = 8'd30;  #10 
a = 8'd104; b = 8'd31;  #10 
a = 8'd104; b = 8'd32;  #10 
a = 8'd104; b = 8'd33;  #10 
a = 8'd104; b = 8'd34;  #10 
a = 8'd104; b = 8'd35;  #10 
a = 8'd104; b = 8'd36;  #10 
a = 8'd104; b = 8'd37;  #10 
a = 8'd104; b = 8'd38;  #10 
a = 8'd104; b = 8'd39;  #10 
a = 8'd104; b = 8'd40;  #10 
a = 8'd104; b = 8'd41;  #10 
a = 8'd104; b = 8'd42;  #10 
a = 8'd104; b = 8'd43;  #10 
a = 8'd104; b = 8'd44;  #10 
a = 8'd104; b = 8'd45;  #10 
a = 8'd104; b = 8'd46;  #10 
a = 8'd104; b = 8'd47;  #10 
a = 8'd104; b = 8'd48;  #10 
a = 8'd104; b = 8'd49;  #10 
a = 8'd104; b = 8'd50;  #10 
a = 8'd104; b = 8'd51;  #10 
a = 8'd104; b = 8'd52;  #10 
a = 8'd104; b = 8'd53;  #10 
a = 8'd104; b = 8'd54;  #10 
a = 8'd104; b = 8'd55;  #10 
a = 8'd104; b = 8'd56;  #10 
a = 8'd104; b = 8'd57;  #10 
a = 8'd104; b = 8'd58;  #10 
a = 8'd104; b = 8'd59;  #10 
a = 8'd104; b = 8'd60;  #10 
a = 8'd104; b = 8'd61;  #10 
a = 8'd104; b = 8'd62;  #10 
a = 8'd104; b = 8'd63;  #10 
a = 8'd104; b = 8'd64;  #10 
a = 8'd104; b = 8'd65;  #10 
a = 8'd104; b = 8'd66;  #10 
a = 8'd104; b = 8'd67;  #10 
a = 8'd104; b = 8'd68;  #10 
a = 8'd104; b = 8'd69;  #10 
a = 8'd104; b = 8'd70;  #10 
a = 8'd104; b = 8'd71;  #10 
a = 8'd104; b = 8'd72;  #10 
a = 8'd104; b = 8'd73;  #10 
a = 8'd104; b = 8'd74;  #10 
a = 8'd104; b = 8'd75;  #10 
a = 8'd104; b = 8'd76;  #10 
a = 8'd104; b = 8'd77;  #10 
a = 8'd104; b = 8'd78;  #10 
a = 8'd104; b = 8'd79;  #10 
a = 8'd104; b = 8'd80;  #10 
a = 8'd104; b = 8'd81;  #10 
a = 8'd104; b = 8'd82;  #10 
a = 8'd104; b = 8'd83;  #10 
a = 8'd104; b = 8'd84;  #10 
a = 8'd104; b = 8'd85;  #10 
a = 8'd104; b = 8'd86;  #10 
a = 8'd104; b = 8'd87;  #10 
a = 8'd104; b = 8'd88;  #10 
a = 8'd104; b = 8'd89;  #10 
a = 8'd104; b = 8'd90;  #10 
a = 8'd104; b = 8'd91;  #10 
a = 8'd104; b = 8'd92;  #10 
a = 8'd104; b = 8'd93;  #10 
a = 8'd104; b = 8'd94;  #10 
a = 8'd104; b = 8'd95;  #10 
a = 8'd104; b = 8'd96;  #10 
a = 8'd104; b = 8'd97;  #10 
a = 8'd104; b = 8'd98;  #10 
a = 8'd104; b = 8'd99;  #10 
a = 8'd104; b = 8'd100;  #10 
a = 8'd104; b = 8'd101;  #10 
a = 8'd104; b = 8'd102;  #10 
a = 8'd104; b = 8'd103;  #10 
a = 8'd104; b = 8'd104;  #10 
a = 8'd104; b = 8'd105;  #10 
a = 8'd104; b = 8'd106;  #10 
a = 8'd104; b = 8'd107;  #10 
a = 8'd104; b = 8'd108;  #10 
a = 8'd104; b = 8'd109;  #10 
a = 8'd104; b = 8'd110;  #10 
a = 8'd104; b = 8'd111;  #10 
a = 8'd104; b = 8'd112;  #10 
a = 8'd104; b = 8'd113;  #10 
a = 8'd104; b = 8'd114;  #10 
a = 8'd104; b = 8'd115;  #10 
a = 8'd104; b = 8'd116;  #10 
a = 8'd104; b = 8'd117;  #10 
a = 8'd104; b = 8'd118;  #10 
a = 8'd104; b = 8'd119;  #10 
a = 8'd104; b = 8'd120;  #10 
a = 8'd104; b = 8'd121;  #10 
a = 8'd104; b = 8'd122;  #10 
a = 8'd104; b = 8'd123;  #10 
a = 8'd104; b = 8'd124;  #10 
a = 8'd104; b = 8'd125;  #10 
a = 8'd104; b = 8'd126;  #10 
a = 8'd104; b = 8'd127;  #10 
a = 8'd104; b = 8'd128;  #10 
a = 8'd104; b = 8'd129;  #10 
a = 8'd104; b = 8'd130;  #10 
a = 8'd104; b = 8'd131;  #10 
a = 8'd104; b = 8'd132;  #10 
a = 8'd104; b = 8'd133;  #10 
a = 8'd104; b = 8'd134;  #10 
a = 8'd104; b = 8'd135;  #10 
a = 8'd104; b = 8'd136;  #10 
a = 8'd104; b = 8'd137;  #10 
a = 8'd104; b = 8'd138;  #10 
a = 8'd104; b = 8'd139;  #10 
a = 8'd104; b = 8'd140;  #10 
a = 8'd104; b = 8'd141;  #10 
a = 8'd104; b = 8'd142;  #10 
a = 8'd104; b = 8'd143;  #10 
a = 8'd104; b = 8'd144;  #10 
a = 8'd104; b = 8'd145;  #10 
a = 8'd104; b = 8'd146;  #10 
a = 8'd104; b = 8'd147;  #10 
a = 8'd104; b = 8'd148;  #10 
a = 8'd104; b = 8'd149;  #10 
a = 8'd104; b = 8'd150;  #10 
a = 8'd104; b = 8'd151;  #10 
a = 8'd104; b = 8'd152;  #10 
a = 8'd104; b = 8'd153;  #10 
a = 8'd104; b = 8'd154;  #10 
a = 8'd104; b = 8'd155;  #10 
a = 8'd104; b = 8'd156;  #10 
a = 8'd104; b = 8'd157;  #10 
a = 8'd104; b = 8'd158;  #10 
a = 8'd104; b = 8'd159;  #10 
a = 8'd104; b = 8'd160;  #10 
a = 8'd104; b = 8'd161;  #10 
a = 8'd104; b = 8'd162;  #10 
a = 8'd104; b = 8'd163;  #10 
a = 8'd104; b = 8'd164;  #10 
a = 8'd104; b = 8'd165;  #10 
a = 8'd104; b = 8'd166;  #10 
a = 8'd104; b = 8'd167;  #10 
a = 8'd104; b = 8'd168;  #10 
a = 8'd104; b = 8'd169;  #10 
a = 8'd104; b = 8'd170;  #10 
a = 8'd104; b = 8'd171;  #10 
a = 8'd104; b = 8'd172;  #10 
a = 8'd104; b = 8'd173;  #10 
a = 8'd104; b = 8'd174;  #10 
a = 8'd104; b = 8'd175;  #10 
a = 8'd104; b = 8'd176;  #10 
a = 8'd104; b = 8'd177;  #10 
a = 8'd104; b = 8'd178;  #10 
a = 8'd104; b = 8'd179;  #10 
a = 8'd104; b = 8'd180;  #10 
a = 8'd104; b = 8'd181;  #10 
a = 8'd104; b = 8'd182;  #10 
a = 8'd104; b = 8'd183;  #10 
a = 8'd104; b = 8'd184;  #10 
a = 8'd104; b = 8'd185;  #10 
a = 8'd104; b = 8'd186;  #10 
a = 8'd104; b = 8'd187;  #10 
a = 8'd104; b = 8'd188;  #10 
a = 8'd104; b = 8'd189;  #10 
a = 8'd104; b = 8'd190;  #10 
a = 8'd104; b = 8'd191;  #10 
a = 8'd104; b = 8'd192;  #10 
a = 8'd104; b = 8'd193;  #10 
a = 8'd104; b = 8'd194;  #10 
a = 8'd104; b = 8'd195;  #10 
a = 8'd104; b = 8'd196;  #10 
a = 8'd104; b = 8'd197;  #10 
a = 8'd104; b = 8'd198;  #10 
a = 8'd104; b = 8'd199;  #10 
a = 8'd104; b = 8'd200;  #10 
a = 8'd104; b = 8'd201;  #10 
a = 8'd104; b = 8'd202;  #10 
a = 8'd104; b = 8'd203;  #10 
a = 8'd104; b = 8'd204;  #10 
a = 8'd104; b = 8'd205;  #10 
a = 8'd104; b = 8'd206;  #10 
a = 8'd104; b = 8'd207;  #10 
a = 8'd104; b = 8'd208;  #10 
a = 8'd104; b = 8'd209;  #10 
a = 8'd104; b = 8'd210;  #10 
a = 8'd104; b = 8'd211;  #10 
a = 8'd104; b = 8'd212;  #10 
a = 8'd104; b = 8'd213;  #10 
a = 8'd104; b = 8'd214;  #10 
a = 8'd104; b = 8'd215;  #10 
a = 8'd104; b = 8'd216;  #10 
a = 8'd104; b = 8'd217;  #10 
a = 8'd104; b = 8'd218;  #10 
a = 8'd104; b = 8'd219;  #10 
a = 8'd104; b = 8'd220;  #10 
a = 8'd104; b = 8'd221;  #10 
a = 8'd104; b = 8'd222;  #10 
a = 8'd104; b = 8'd223;  #10 
a = 8'd104; b = 8'd224;  #10 
a = 8'd104; b = 8'd225;  #10 
a = 8'd104; b = 8'd226;  #10 
a = 8'd104; b = 8'd227;  #10 
a = 8'd104; b = 8'd228;  #10 
a = 8'd104; b = 8'd229;  #10 
a = 8'd104; b = 8'd230;  #10 
a = 8'd104; b = 8'd231;  #10 
a = 8'd104; b = 8'd232;  #10 
a = 8'd104; b = 8'd233;  #10 
a = 8'd104; b = 8'd234;  #10 
a = 8'd104; b = 8'd235;  #10 
a = 8'd104; b = 8'd236;  #10 
a = 8'd104; b = 8'd237;  #10 
a = 8'd104; b = 8'd238;  #10 
a = 8'd104; b = 8'd239;  #10 
a = 8'd104; b = 8'd240;  #10 
a = 8'd104; b = 8'd241;  #10 
a = 8'd104; b = 8'd242;  #10 
a = 8'd104; b = 8'd243;  #10 
a = 8'd104; b = 8'd244;  #10 
a = 8'd104; b = 8'd245;  #10 
a = 8'd104; b = 8'd246;  #10 
a = 8'd104; b = 8'd247;  #10 
a = 8'd104; b = 8'd248;  #10 
a = 8'd104; b = 8'd249;  #10 
a = 8'd104; b = 8'd250;  #10 
a = 8'd104; b = 8'd251;  #10 
a = 8'd104; b = 8'd252;  #10 
a = 8'd104; b = 8'd253;  #10 
a = 8'd104; b = 8'd254;  #10 
a = 8'd104; b = 8'd255;  #10 
a = 8'd105; b = 8'd0;  #10 
a = 8'd105; b = 8'd1;  #10 
a = 8'd105; b = 8'd2;  #10 
a = 8'd105; b = 8'd3;  #10 
a = 8'd105; b = 8'd4;  #10 
a = 8'd105; b = 8'd5;  #10 
a = 8'd105; b = 8'd6;  #10 
a = 8'd105; b = 8'd7;  #10 
a = 8'd105; b = 8'd8;  #10 
a = 8'd105; b = 8'd9;  #10 
a = 8'd105; b = 8'd10;  #10 
a = 8'd105; b = 8'd11;  #10 
a = 8'd105; b = 8'd12;  #10 
a = 8'd105; b = 8'd13;  #10 
a = 8'd105; b = 8'd14;  #10 
a = 8'd105; b = 8'd15;  #10 
a = 8'd105; b = 8'd16;  #10 
a = 8'd105; b = 8'd17;  #10 
a = 8'd105; b = 8'd18;  #10 
a = 8'd105; b = 8'd19;  #10 
a = 8'd105; b = 8'd20;  #10 
a = 8'd105; b = 8'd21;  #10 
a = 8'd105; b = 8'd22;  #10 
a = 8'd105; b = 8'd23;  #10 
a = 8'd105; b = 8'd24;  #10 
a = 8'd105; b = 8'd25;  #10 
a = 8'd105; b = 8'd26;  #10 
a = 8'd105; b = 8'd27;  #10 
a = 8'd105; b = 8'd28;  #10 
a = 8'd105; b = 8'd29;  #10 
a = 8'd105; b = 8'd30;  #10 
a = 8'd105; b = 8'd31;  #10 
a = 8'd105; b = 8'd32;  #10 
a = 8'd105; b = 8'd33;  #10 
a = 8'd105; b = 8'd34;  #10 
a = 8'd105; b = 8'd35;  #10 
a = 8'd105; b = 8'd36;  #10 
a = 8'd105; b = 8'd37;  #10 
a = 8'd105; b = 8'd38;  #10 
a = 8'd105; b = 8'd39;  #10 
a = 8'd105; b = 8'd40;  #10 
a = 8'd105; b = 8'd41;  #10 
a = 8'd105; b = 8'd42;  #10 
a = 8'd105; b = 8'd43;  #10 
a = 8'd105; b = 8'd44;  #10 
a = 8'd105; b = 8'd45;  #10 
a = 8'd105; b = 8'd46;  #10 
a = 8'd105; b = 8'd47;  #10 
a = 8'd105; b = 8'd48;  #10 
a = 8'd105; b = 8'd49;  #10 
a = 8'd105; b = 8'd50;  #10 
a = 8'd105; b = 8'd51;  #10 
a = 8'd105; b = 8'd52;  #10 
a = 8'd105; b = 8'd53;  #10 
a = 8'd105; b = 8'd54;  #10 
a = 8'd105; b = 8'd55;  #10 
a = 8'd105; b = 8'd56;  #10 
a = 8'd105; b = 8'd57;  #10 
a = 8'd105; b = 8'd58;  #10 
a = 8'd105; b = 8'd59;  #10 
a = 8'd105; b = 8'd60;  #10 
a = 8'd105; b = 8'd61;  #10 
a = 8'd105; b = 8'd62;  #10 
a = 8'd105; b = 8'd63;  #10 
a = 8'd105; b = 8'd64;  #10 
a = 8'd105; b = 8'd65;  #10 
a = 8'd105; b = 8'd66;  #10 
a = 8'd105; b = 8'd67;  #10 
a = 8'd105; b = 8'd68;  #10 
a = 8'd105; b = 8'd69;  #10 
a = 8'd105; b = 8'd70;  #10 
a = 8'd105; b = 8'd71;  #10 
a = 8'd105; b = 8'd72;  #10 
a = 8'd105; b = 8'd73;  #10 
a = 8'd105; b = 8'd74;  #10 
a = 8'd105; b = 8'd75;  #10 
a = 8'd105; b = 8'd76;  #10 
a = 8'd105; b = 8'd77;  #10 
a = 8'd105; b = 8'd78;  #10 
a = 8'd105; b = 8'd79;  #10 
a = 8'd105; b = 8'd80;  #10 
a = 8'd105; b = 8'd81;  #10 
a = 8'd105; b = 8'd82;  #10 
a = 8'd105; b = 8'd83;  #10 
a = 8'd105; b = 8'd84;  #10 
a = 8'd105; b = 8'd85;  #10 
a = 8'd105; b = 8'd86;  #10 
a = 8'd105; b = 8'd87;  #10 
a = 8'd105; b = 8'd88;  #10 
a = 8'd105; b = 8'd89;  #10 
a = 8'd105; b = 8'd90;  #10 
a = 8'd105; b = 8'd91;  #10 
a = 8'd105; b = 8'd92;  #10 
a = 8'd105; b = 8'd93;  #10 
a = 8'd105; b = 8'd94;  #10 
a = 8'd105; b = 8'd95;  #10 
a = 8'd105; b = 8'd96;  #10 
a = 8'd105; b = 8'd97;  #10 
a = 8'd105; b = 8'd98;  #10 
a = 8'd105; b = 8'd99;  #10 
a = 8'd105; b = 8'd100;  #10 
a = 8'd105; b = 8'd101;  #10 
a = 8'd105; b = 8'd102;  #10 
a = 8'd105; b = 8'd103;  #10 
a = 8'd105; b = 8'd104;  #10 
a = 8'd105; b = 8'd105;  #10 
a = 8'd105; b = 8'd106;  #10 
a = 8'd105; b = 8'd107;  #10 
a = 8'd105; b = 8'd108;  #10 
a = 8'd105; b = 8'd109;  #10 
a = 8'd105; b = 8'd110;  #10 
a = 8'd105; b = 8'd111;  #10 
a = 8'd105; b = 8'd112;  #10 
a = 8'd105; b = 8'd113;  #10 
a = 8'd105; b = 8'd114;  #10 
a = 8'd105; b = 8'd115;  #10 
a = 8'd105; b = 8'd116;  #10 
a = 8'd105; b = 8'd117;  #10 
a = 8'd105; b = 8'd118;  #10 
a = 8'd105; b = 8'd119;  #10 
a = 8'd105; b = 8'd120;  #10 
a = 8'd105; b = 8'd121;  #10 
a = 8'd105; b = 8'd122;  #10 
a = 8'd105; b = 8'd123;  #10 
a = 8'd105; b = 8'd124;  #10 
a = 8'd105; b = 8'd125;  #10 
a = 8'd105; b = 8'd126;  #10 
a = 8'd105; b = 8'd127;  #10 
a = 8'd105; b = 8'd128;  #10 
a = 8'd105; b = 8'd129;  #10 
a = 8'd105; b = 8'd130;  #10 
a = 8'd105; b = 8'd131;  #10 
a = 8'd105; b = 8'd132;  #10 
a = 8'd105; b = 8'd133;  #10 
a = 8'd105; b = 8'd134;  #10 
a = 8'd105; b = 8'd135;  #10 
a = 8'd105; b = 8'd136;  #10 
a = 8'd105; b = 8'd137;  #10 
a = 8'd105; b = 8'd138;  #10 
a = 8'd105; b = 8'd139;  #10 
a = 8'd105; b = 8'd140;  #10 
a = 8'd105; b = 8'd141;  #10 
a = 8'd105; b = 8'd142;  #10 
a = 8'd105; b = 8'd143;  #10 
a = 8'd105; b = 8'd144;  #10 
a = 8'd105; b = 8'd145;  #10 
a = 8'd105; b = 8'd146;  #10 
a = 8'd105; b = 8'd147;  #10 
a = 8'd105; b = 8'd148;  #10 
a = 8'd105; b = 8'd149;  #10 
a = 8'd105; b = 8'd150;  #10 
a = 8'd105; b = 8'd151;  #10 
a = 8'd105; b = 8'd152;  #10 
a = 8'd105; b = 8'd153;  #10 
a = 8'd105; b = 8'd154;  #10 
a = 8'd105; b = 8'd155;  #10 
a = 8'd105; b = 8'd156;  #10 
a = 8'd105; b = 8'd157;  #10 
a = 8'd105; b = 8'd158;  #10 
a = 8'd105; b = 8'd159;  #10 
a = 8'd105; b = 8'd160;  #10 
a = 8'd105; b = 8'd161;  #10 
a = 8'd105; b = 8'd162;  #10 
a = 8'd105; b = 8'd163;  #10 
a = 8'd105; b = 8'd164;  #10 
a = 8'd105; b = 8'd165;  #10 
a = 8'd105; b = 8'd166;  #10 
a = 8'd105; b = 8'd167;  #10 
a = 8'd105; b = 8'd168;  #10 
a = 8'd105; b = 8'd169;  #10 
a = 8'd105; b = 8'd170;  #10 
a = 8'd105; b = 8'd171;  #10 
a = 8'd105; b = 8'd172;  #10 
a = 8'd105; b = 8'd173;  #10 
a = 8'd105; b = 8'd174;  #10 
a = 8'd105; b = 8'd175;  #10 
a = 8'd105; b = 8'd176;  #10 
a = 8'd105; b = 8'd177;  #10 
a = 8'd105; b = 8'd178;  #10 
a = 8'd105; b = 8'd179;  #10 
a = 8'd105; b = 8'd180;  #10 
a = 8'd105; b = 8'd181;  #10 
a = 8'd105; b = 8'd182;  #10 
a = 8'd105; b = 8'd183;  #10 
a = 8'd105; b = 8'd184;  #10 
a = 8'd105; b = 8'd185;  #10 
a = 8'd105; b = 8'd186;  #10 
a = 8'd105; b = 8'd187;  #10 
a = 8'd105; b = 8'd188;  #10 
a = 8'd105; b = 8'd189;  #10 
a = 8'd105; b = 8'd190;  #10 
a = 8'd105; b = 8'd191;  #10 
a = 8'd105; b = 8'd192;  #10 
a = 8'd105; b = 8'd193;  #10 
a = 8'd105; b = 8'd194;  #10 
a = 8'd105; b = 8'd195;  #10 
a = 8'd105; b = 8'd196;  #10 
a = 8'd105; b = 8'd197;  #10 
a = 8'd105; b = 8'd198;  #10 
a = 8'd105; b = 8'd199;  #10 
a = 8'd105; b = 8'd200;  #10 
a = 8'd105; b = 8'd201;  #10 
a = 8'd105; b = 8'd202;  #10 
a = 8'd105; b = 8'd203;  #10 
a = 8'd105; b = 8'd204;  #10 
a = 8'd105; b = 8'd205;  #10 
a = 8'd105; b = 8'd206;  #10 
a = 8'd105; b = 8'd207;  #10 
a = 8'd105; b = 8'd208;  #10 
a = 8'd105; b = 8'd209;  #10 
a = 8'd105; b = 8'd210;  #10 
a = 8'd105; b = 8'd211;  #10 
a = 8'd105; b = 8'd212;  #10 
a = 8'd105; b = 8'd213;  #10 
a = 8'd105; b = 8'd214;  #10 
a = 8'd105; b = 8'd215;  #10 
a = 8'd105; b = 8'd216;  #10 
a = 8'd105; b = 8'd217;  #10 
a = 8'd105; b = 8'd218;  #10 
a = 8'd105; b = 8'd219;  #10 
a = 8'd105; b = 8'd220;  #10 
a = 8'd105; b = 8'd221;  #10 
a = 8'd105; b = 8'd222;  #10 
a = 8'd105; b = 8'd223;  #10 
a = 8'd105; b = 8'd224;  #10 
a = 8'd105; b = 8'd225;  #10 
a = 8'd105; b = 8'd226;  #10 
a = 8'd105; b = 8'd227;  #10 
a = 8'd105; b = 8'd228;  #10 
a = 8'd105; b = 8'd229;  #10 
a = 8'd105; b = 8'd230;  #10 
a = 8'd105; b = 8'd231;  #10 
a = 8'd105; b = 8'd232;  #10 
a = 8'd105; b = 8'd233;  #10 
a = 8'd105; b = 8'd234;  #10 
a = 8'd105; b = 8'd235;  #10 
a = 8'd105; b = 8'd236;  #10 
a = 8'd105; b = 8'd237;  #10 
a = 8'd105; b = 8'd238;  #10 
a = 8'd105; b = 8'd239;  #10 
a = 8'd105; b = 8'd240;  #10 
a = 8'd105; b = 8'd241;  #10 
a = 8'd105; b = 8'd242;  #10 
a = 8'd105; b = 8'd243;  #10 
a = 8'd105; b = 8'd244;  #10 
a = 8'd105; b = 8'd245;  #10 
a = 8'd105; b = 8'd246;  #10 
a = 8'd105; b = 8'd247;  #10 
a = 8'd105; b = 8'd248;  #10 
a = 8'd105; b = 8'd249;  #10 
a = 8'd105; b = 8'd250;  #10 
a = 8'd105; b = 8'd251;  #10 
a = 8'd105; b = 8'd252;  #10 
a = 8'd105; b = 8'd253;  #10 
a = 8'd105; b = 8'd254;  #10 
a = 8'd105; b = 8'd255;  #10 
a = 8'd106; b = 8'd0;  #10 
a = 8'd106; b = 8'd1;  #10 
a = 8'd106; b = 8'd2;  #10 
a = 8'd106; b = 8'd3;  #10 
a = 8'd106; b = 8'd4;  #10 
a = 8'd106; b = 8'd5;  #10 
a = 8'd106; b = 8'd6;  #10 
a = 8'd106; b = 8'd7;  #10 
a = 8'd106; b = 8'd8;  #10 
a = 8'd106; b = 8'd9;  #10 
a = 8'd106; b = 8'd10;  #10 
a = 8'd106; b = 8'd11;  #10 
a = 8'd106; b = 8'd12;  #10 
a = 8'd106; b = 8'd13;  #10 
a = 8'd106; b = 8'd14;  #10 
a = 8'd106; b = 8'd15;  #10 
a = 8'd106; b = 8'd16;  #10 
a = 8'd106; b = 8'd17;  #10 
a = 8'd106; b = 8'd18;  #10 
a = 8'd106; b = 8'd19;  #10 
a = 8'd106; b = 8'd20;  #10 
a = 8'd106; b = 8'd21;  #10 
a = 8'd106; b = 8'd22;  #10 
a = 8'd106; b = 8'd23;  #10 
a = 8'd106; b = 8'd24;  #10 
a = 8'd106; b = 8'd25;  #10 
a = 8'd106; b = 8'd26;  #10 
a = 8'd106; b = 8'd27;  #10 
a = 8'd106; b = 8'd28;  #10 
a = 8'd106; b = 8'd29;  #10 
a = 8'd106; b = 8'd30;  #10 
a = 8'd106; b = 8'd31;  #10 
a = 8'd106; b = 8'd32;  #10 
a = 8'd106; b = 8'd33;  #10 
a = 8'd106; b = 8'd34;  #10 
a = 8'd106; b = 8'd35;  #10 
a = 8'd106; b = 8'd36;  #10 
a = 8'd106; b = 8'd37;  #10 
a = 8'd106; b = 8'd38;  #10 
a = 8'd106; b = 8'd39;  #10 
a = 8'd106; b = 8'd40;  #10 
a = 8'd106; b = 8'd41;  #10 
a = 8'd106; b = 8'd42;  #10 
a = 8'd106; b = 8'd43;  #10 
a = 8'd106; b = 8'd44;  #10 
a = 8'd106; b = 8'd45;  #10 
a = 8'd106; b = 8'd46;  #10 
a = 8'd106; b = 8'd47;  #10 
a = 8'd106; b = 8'd48;  #10 
a = 8'd106; b = 8'd49;  #10 
a = 8'd106; b = 8'd50;  #10 
a = 8'd106; b = 8'd51;  #10 
a = 8'd106; b = 8'd52;  #10 
a = 8'd106; b = 8'd53;  #10 
a = 8'd106; b = 8'd54;  #10 
a = 8'd106; b = 8'd55;  #10 
a = 8'd106; b = 8'd56;  #10 
a = 8'd106; b = 8'd57;  #10 
a = 8'd106; b = 8'd58;  #10 
a = 8'd106; b = 8'd59;  #10 
a = 8'd106; b = 8'd60;  #10 
a = 8'd106; b = 8'd61;  #10 
a = 8'd106; b = 8'd62;  #10 
a = 8'd106; b = 8'd63;  #10 
a = 8'd106; b = 8'd64;  #10 
a = 8'd106; b = 8'd65;  #10 
a = 8'd106; b = 8'd66;  #10 
a = 8'd106; b = 8'd67;  #10 
a = 8'd106; b = 8'd68;  #10 
a = 8'd106; b = 8'd69;  #10 
a = 8'd106; b = 8'd70;  #10 
a = 8'd106; b = 8'd71;  #10 
a = 8'd106; b = 8'd72;  #10 
a = 8'd106; b = 8'd73;  #10 
a = 8'd106; b = 8'd74;  #10 
a = 8'd106; b = 8'd75;  #10 
a = 8'd106; b = 8'd76;  #10 
a = 8'd106; b = 8'd77;  #10 
a = 8'd106; b = 8'd78;  #10 
a = 8'd106; b = 8'd79;  #10 
a = 8'd106; b = 8'd80;  #10 
a = 8'd106; b = 8'd81;  #10 
a = 8'd106; b = 8'd82;  #10 
a = 8'd106; b = 8'd83;  #10 
a = 8'd106; b = 8'd84;  #10 
a = 8'd106; b = 8'd85;  #10 
a = 8'd106; b = 8'd86;  #10 
a = 8'd106; b = 8'd87;  #10 
a = 8'd106; b = 8'd88;  #10 
a = 8'd106; b = 8'd89;  #10 
a = 8'd106; b = 8'd90;  #10 
a = 8'd106; b = 8'd91;  #10 
a = 8'd106; b = 8'd92;  #10 
a = 8'd106; b = 8'd93;  #10 
a = 8'd106; b = 8'd94;  #10 
a = 8'd106; b = 8'd95;  #10 
a = 8'd106; b = 8'd96;  #10 
a = 8'd106; b = 8'd97;  #10 
a = 8'd106; b = 8'd98;  #10 
a = 8'd106; b = 8'd99;  #10 
a = 8'd106; b = 8'd100;  #10 
a = 8'd106; b = 8'd101;  #10 
a = 8'd106; b = 8'd102;  #10 
a = 8'd106; b = 8'd103;  #10 
a = 8'd106; b = 8'd104;  #10 
a = 8'd106; b = 8'd105;  #10 
a = 8'd106; b = 8'd106;  #10 
a = 8'd106; b = 8'd107;  #10 
a = 8'd106; b = 8'd108;  #10 
a = 8'd106; b = 8'd109;  #10 
a = 8'd106; b = 8'd110;  #10 
a = 8'd106; b = 8'd111;  #10 
a = 8'd106; b = 8'd112;  #10 
a = 8'd106; b = 8'd113;  #10 
a = 8'd106; b = 8'd114;  #10 
a = 8'd106; b = 8'd115;  #10 
a = 8'd106; b = 8'd116;  #10 
a = 8'd106; b = 8'd117;  #10 
a = 8'd106; b = 8'd118;  #10 
a = 8'd106; b = 8'd119;  #10 
a = 8'd106; b = 8'd120;  #10 
a = 8'd106; b = 8'd121;  #10 
a = 8'd106; b = 8'd122;  #10 
a = 8'd106; b = 8'd123;  #10 
a = 8'd106; b = 8'd124;  #10 
a = 8'd106; b = 8'd125;  #10 
a = 8'd106; b = 8'd126;  #10 
a = 8'd106; b = 8'd127;  #10 
a = 8'd106; b = 8'd128;  #10 
a = 8'd106; b = 8'd129;  #10 
a = 8'd106; b = 8'd130;  #10 
a = 8'd106; b = 8'd131;  #10 
a = 8'd106; b = 8'd132;  #10 
a = 8'd106; b = 8'd133;  #10 
a = 8'd106; b = 8'd134;  #10 
a = 8'd106; b = 8'd135;  #10 
a = 8'd106; b = 8'd136;  #10 
a = 8'd106; b = 8'd137;  #10 
a = 8'd106; b = 8'd138;  #10 
a = 8'd106; b = 8'd139;  #10 
a = 8'd106; b = 8'd140;  #10 
a = 8'd106; b = 8'd141;  #10 
a = 8'd106; b = 8'd142;  #10 
a = 8'd106; b = 8'd143;  #10 
a = 8'd106; b = 8'd144;  #10 
a = 8'd106; b = 8'd145;  #10 
a = 8'd106; b = 8'd146;  #10 
a = 8'd106; b = 8'd147;  #10 
a = 8'd106; b = 8'd148;  #10 
a = 8'd106; b = 8'd149;  #10 
a = 8'd106; b = 8'd150;  #10 
a = 8'd106; b = 8'd151;  #10 
a = 8'd106; b = 8'd152;  #10 
a = 8'd106; b = 8'd153;  #10 
a = 8'd106; b = 8'd154;  #10 
a = 8'd106; b = 8'd155;  #10 
a = 8'd106; b = 8'd156;  #10 
a = 8'd106; b = 8'd157;  #10 
a = 8'd106; b = 8'd158;  #10 
a = 8'd106; b = 8'd159;  #10 
a = 8'd106; b = 8'd160;  #10 
a = 8'd106; b = 8'd161;  #10 
a = 8'd106; b = 8'd162;  #10 
a = 8'd106; b = 8'd163;  #10 
a = 8'd106; b = 8'd164;  #10 
a = 8'd106; b = 8'd165;  #10 
a = 8'd106; b = 8'd166;  #10 
a = 8'd106; b = 8'd167;  #10 
a = 8'd106; b = 8'd168;  #10 
a = 8'd106; b = 8'd169;  #10 
a = 8'd106; b = 8'd170;  #10 
a = 8'd106; b = 8'd171;  #10 
a = 8'd106; b = 8'd172;  #10 
a = 8'd106; b = 8'd173;  #10 
a = 8'd106; b = 8'd174;  #10 
a = 8'd106; b = 8'd175;  #10 
a = 8'd106; b = 8'd176;  #10 
a = 8'd106; b = 8'd177;  #10 
a = 8'd106; b = 8'd178;  #10 
a = 8'd106; b = 8'd179;  #10 
a = 8'd106; b = 8'd180;  #10 
a = 8'd106; b = 8'd181;  #10 
a = 8'd106; b = 8'd182;  #10 
a = 8'd106; b = 8'd183;  #10 
a = 8'd106; b = 8'd184;  #10 
a = 8'd106; b = 8'd185;  #10 
a = 8'd106; b = 8'd186;  #10 
a = 8'd106; b = 8'd187;  #10 
a = 8'd106; b = 8'd188;  #10 
a = 8'd106; b = 8'd189;  #10 
a = 8'd106; b = 8'd190;  #10 
a = 8'd106; b = 8'd191;  #10 
a = 8'd106; b = 8'd192;  #10 
a = 8'd106; b = 8'd193;  #10 
a = 8'd106; b = 8'd194;  #10 
a = 8'd106; b = 8'd195;  #10 
a = 8'd106; b = 8'd196;  #10 
a = 8'd106; b = 8'd197;  #10 
a = 8'd106; b = 8'd198;  #10 
a = 8'd106; b = 8'd199;  #10 
a = 8'd106; b = 8'd200;  #10 
a = 8'd106; b = 8'd201;  #10 
a = 8'd106; b = 8'd202;  #10 
a = 8'd106; b = 8'd203;  #10 
a = 8'd106; b = 8'd204;  #10 
a = 8'd106; b = 8'd205;  #10 
a = 8'd106; b = 8'd206;  #10 
a = 8'd106; b = 8'd207;  #10 
a = 8'd106; b = 8'd208;  #10 
a = 8'd106; b = 8'd209;  #10 
a = 8'd106; b = 8'd210;  #10 
a = 8'd106; b = 8'd211;  #10 
a = 8'd106; b = 8'd212;  #10 
a = 8'd106; b = 8'd213;  #10 
a = 8'd106; b = 8'd214;  #10 
a = 8'd106; b = 8'd215;  #10 
a = 8'd106; b = 8'd216;  #10 
a = 8'd106; b = 8'd217;  #10 
a = 8'd106; b = 8'd218;  #10 
a = 8'd106; b = 8'd219;  #10 
a = 8'd106; b = 8'd220;  #10 
a = 8'd106; b = 8'd221;  #10 
a = 8'd106; b = 8'd222;  #10 
a = 8'd106; b = 8'd223;  #10 
a = 8'd106; b = 8'd224;  #10 
a = 8'd106; b = 8'd225;  #10 
a = 8'd106; b = 8'd226;  #10 
a = 8'd106; b = 8'd227;  #10 
a = 8'd106; b = 8'd228;  #10 
a = 8'd106; b = 8'd229;  #10 
a = 8'd106; b = 8'd230;  #10 
a = 8'd106; b = 8'd231;  #10 
a = 8'd106; b = 8'd232;  #10 
a = 8'd106; b = 8'd233;  #10 
a = 8'd106; b = 8'd234;  #10 
a = 8'd106; b = 8'd235;  #10 
a = 8'd106; b = 8'd236;  #10 
a = 8'd106; b = 8'd237;  #10 
a = 8'd106; b = 8'd238;  #10 
a = 8'd106; b = 8'd239;  #10 
a = 8'd106; b = 8'd240;  #10 
a = 8'd106; b = 8'd241;  #10 
a = 8'd106; b = 8'd242;  #10 
a = 8'd106; b = 8'd243;  #10 
a = 8'd106; b = 8'd244;  #10 
a = 8'd106; b = 8'd245;  #10 
a = 8'd106; b = 8'd246;  #10 
a = 8'd106; b = 8'd247;  #10 
a = 8'd106; b = 8'd248;  #10 
a = 8'd106; b = 8'd249;  #10 
a = 8'd106; b = 8'd250;  #10 
a = 8'd106; b = 8'd251;  #10 
a = 8'd106; b = 8'd252;  #10 
a = 8'd106; b = 8'd253;  #10 
a = 8'd106; b = 8'd254;  #10 
a = 8'd106; b = 8'd255;  #10 
a = 8'd107; b = 8'd0;  #10 
a = 8'd107; b = 8'd1;  #10 
a = 8'd107; b = 8'd2;  #10 
a = 8'd107; b = 8'd3;  #10 
a = 8'd107; b = 8'd4;  #10 
a = 8'd107; b = 8'd5;  #10 
a = 8'd107; b = 8'd6;  #10 
a = 8'd107; b = 8'd7;  #10 
a = 8'd107; b = 8'd8;  #10 
a = 8'd107; b = 8'd9;  #10 
a = 8'd107; b = 8'd10;  #10 
a = 8'd107; b = 8'd11;  #10 
a = 8'd107; b = 8'd12;  #10 
a = 8'd107; b = 8'd13;  #10 
a = 8'd107; b = 8'd14;  #10 
a = 8'd107; b = 8'd15;  #10 
a = 8'd107; b = 8'd16;  #10 
a = 8'd107; b = 8'd17;  #10 
a = 8'd107; b = 8'd18;  #10 
a = 8'd107; b = 8'd19;  #10 
a = 8'd107; b = 8'd20;  #10 
a = 8'd107; b = 8'd21;  #10 
a = 8'd107; b = 8'd22;  #10 
a = 8'd107; b = 8'd23;  #10 
a = 8'd107; b = 8'd24;  #10 
a = 8'd107; b = 8'd25;  #10 
a = 8'd107; b = 8'd26;  #10 
a = 8'd107; b = 8'd27;  #10 
a = 8'd107; b = 8'd28;  #10 
a = 8'd107; b = 8'd29;  #10 
a = 8'd107; b = 8'd30;  #10 
a = 8'd107; b = 8'd31;  #10 
a = 8'd107; b = 8'd32;  #10 
a = 8'd107; b = 8'd33;  #10 
a = 8'd107; b = 8'd34;  #10 
a = 8'd107; b = 8'd35;  #10 
a = 8'd107; b = 8'd36;  #10 
a = 8'd107; b = 8'd37;  #10 
a = 8'd107; b = 8'd38;  #10 
a = 8'd107; b = 8'd39;  #10 
a = 8'd107; b = 8'd40;  #10 
a = 8'd107; b = 8'd41;  #10 
a = 8'd107; b = 8'd42;  #10 
a = 8'd107; b = 8'd43;  #10 
a = 8'd107; b = 8'd44;  #10 
a = 8'd107; b = 8'd45;  #10 
a = 8'd107; b = 8'd46;  #10 
a = 8'd107; b = 8'd47;  #10 
a = 8'd107; b = 8'd48;  #10 
a = 8'd107; b = 8'd49;  #10 
a = 8'd107; b = 8'd50;  #10 
a = 8'd107; b = 8'd51;  #10 
a = 8'd107; b = 8'd52;  #10 
a = 8'd107; b = 8'd53;  #10 
a = 8'd107; b = 8'd54;  #10 
a = 8'd107; b = 8'd55;  #10 
a = 8'd107; b = 8'd56;  #10 
a = 8'd107; b = 8'd57;  #10 
a = 8'd107; b = 8'd58;  #10 
a = 8'd107; b = 8'd59;  #10 
a = 8'd107; b = 8'd60;  #10 
a = 8'd107; b = 8'd61;  #10 
a = 8'd107; b = 8'd62;  #10 
a = 8'd107; b = 8'd63;  #10 
a = 8'd107; b = 8'd64;  #10 
a = 8'd107; b = 8'd65;  #10 
a = 8'd107; b = 8'd66;  #10 
a = 8'd107; b = 8'd67;  #10 
a = 8'd107; b = 8'd68;  #10 
a = 8'd107; b = 8'd69;  #10 
a = 8'd107; b = 8'd70;  #10 
a = 8'd107; b = 8'd71;  #10 
a = 8'd107; b = 8'd72;  #10 
a = 8'd107; b = 8'd73;  #10 
a = 8'd107; b = 8'd74;  #10 
a = 8'd107; b = 8'd75;  #10 
a = 8'd107; b = 8'd76;  #10 
a = 8'd107; b = 8'd77;  #10 
a = 8'd107; b = 8'd78;  #10 
a = 8'd107; b = 8'd79;  #10 
a = 8'd107; b = 8'd80;  #10 
a = 8'd107; b = 8'd81;  #10 
a = 8'd107; b = 8'd82;  #10 
a = 8'd107; b = 8'd83;  #10 
a = 8'd107; b = 8'd84;  #10 
a = 8'd107; b = 8'd85;  #10 
a = 8'd107; b = 8'd86;  #10 
a = 8'd107; b = 8'd87;  #10 
a = 8'd107; b = 8'd88;  #10 
a = 8'd107; b = 8'd89;  #10 
a = 8'd107; b = 8'd90;  #10 
a = 8'd107; b = 8'd91;  #10 
a = 8'd107; b = 8'd92;  #10 
a = 8'd107; b = 8'd93;  #10 
a = 8'd107; b = 8'd94;  #10 
a = 8'd107; b = 8'd95;  #10 
a = 8'd107; b = 8'd96;  #10 
a = 8'd107; b = 8'd97;  #10 
a = 8'd107; b = 8'd98;  #10 
a = 8'd107; b = 8'd99;  #10 
a = 8'd107; b = 8'd100;  #10 
a = 8'd107; b = 8'd101;  #10 
a = 8'd107; b = 8'd102;  #10 
a = 8'd107; b = 8'd103;  #10 
a = 8'd107; b = 8'd104;  #10 
a = 8'd107; b = 8'd105;  #10 
a = 8'd107; b = 8'd106;  #10 
a = 8'd107; b = 8'd107;  #10 
a = 8'd107; b = 8'd108;  #10 
a = 8'd107; b = 8'd109;  #10 
a = 8'd107; b = 8'd110;  #10 
a = 8'd107; b = 8'd111;  #10 
a = 8'd107; b = 8'd112;  #10 
a = 8'd107; b = 8'd113;  #10 
a = 8'd107; b = 8'd114;  #10 
a = 8'd107; b = 8'd115;  #10 
a = 8'd107; b = 8'd116;  #10 
a = 8'd107; b = 8'd117;  #10 
a = 8'd107; b = 8'd118;  #10 
a = 8'd107; b = 8'd119;  #10 
a = 8'd107; b = 8'd120;  #10 
a = 8'd107; b = 8'd121;  #10 
a = 8'd107; b = 8'd122;  #10 
a = 8'd107; b = 8'd123;  #10 
a = 8'd107; b = 8'd124;  #10 
a = 8'd107; b = 8'd125;  #10 
a = 8'd107; b = 8'd126;  #10 
a = 8'd107; b = 8'd127;  #10 
a = 8'd107; b = 8'd128;  #10 
a = 8'd107; b = 8'd129;  #10 
a = 8'd107; b = 8'd130;  #10 
a = 8'd107; b = 8'd131;  #10 
a = 8'd107; b = 8'd132;  #10 
a = 8'd107; b = 8'd133;  #10 
a = 8'd107; b = 8'd134;  #10 
a = 8'd107; b = 8'd135;  #10 
a = 8'd107; b = 8'd136;  #10 
a = 8'd107; b = 8'd137;  #10 
a = 8'd107; b = 8'd138;  #10 
a = 8'd107; b = 8'd139;  #10 
a = 8'd107; b = 8'd140;  #10 
a = 8'd107; b = 8'd141;  #10 
a = 8'd107; b = 8'd142;  #10 
a = 8'd107; b = 8'd143;  #10 
a = 8'd107; b = 8'd144;  #10 
a = 8'd107; b = 8'd145;  #10 
a = 8'd107; b = 8'd146;  #10 
a = 8'd107; b = 8'd147;  #10 
a = 8'd107; b = 8'd148;  #10 
a = 8'd107; b = 8'd149;  #10 
a = 8'd107; b = 8'd150;  #10 
a = 8'd107; b = 8'd151;  #10 
a = 8'd107; b = 8'd152;  #10 
a = 8'd107; b = 8'd153;  #10 
a = 8'd107; b = 8'd154;  #10 
a = 8'd107; b = 8'd155;  #10 
a = 8'd107; b = 8'd156;  #10 
a = 8'd107; b = 8'd157;  #10 
a = 8'd107; b = 8'd158;  #10 
a = 8'd107; b = 8'd159;  #10 
a = 8'd107; b = 8'd160;  #10 
a = 8'd107; b = 8'd161;  #10 
a = 8'd107; b = 8'd162;  #10 
a = 8'd107; b = 8'd163;  #10 
a = 8'd107; b = 8'd164;  #10 
a = 8'd107; b = 8'd165;  #10 
a = 8'd107; b = 8'd166;  #10 
a = 8'd107; b = 8'd167;  #10 
a = 8'd107; b = 8'd168;  #10 
a = 8'd107; b = 8'd169;  #10 
a = 8'd107; b = 8'd170;  #10 
a = 8'd107; b = 8'd171;  #10 
a = 8'd107; b = 8'd172;  #10 
a = 8'd107; b = 8'd173;  #10 
a = 8'd107; b = 8'd174;  #10 
a = 8'd107; b = 8'd175;  #10 
a = 8'd107; b = 8'd176;  #10 
a = 8'd107; b = 8'd177;  #10 
a = 8'd107; b = 8'd178;  #10 
a = 8'd107; b = 8'd179;  #10 
a = 8'd107; b = 8'd180;  #10 
a = 8'd107; b = 8'd181;  #10 
a = 8'd107; b = 8'd182;  #10 
a = 8'd107; b = 8'd183;  #10 
a = 8'd107; b = 8'd184;  #10 
a = 8'd107; b = 8'd185;  #10 
a = 8'd107; b = 8'd186;  #10 
a = 8'd107; b = 8'd187;  #10 
a = 8'd107; b = 8'd188;  #10 
a = 8'd107; b = 8'd189;  #10 
a = 8'd107; b = 8'd190;  #10 
a = 8'd107; b = 8'd191;  #10 
a = 8'd107; b = 8'd192;  #10 
a = 8'd107; b = 8'd193;  #10 
a = 8'd107; b = 8'd194;  #10 
a = 8'd107; b = 8'd195;  #10 
a = 8'd107; b = 8'd196;  #10 
a = 8'd107; b = 8'd197;  #10 
a = 8'd107; b = 8'd198;  #10 
a = 8'd107; b = 8'd199;  #10 
a = 8'd107; b = 8'd200;  #10 
a = 8'd107; b = 8'd201;  #10 
a = 8'd107; b = 8'd202;  #10 
a = 8'd107; b = 8'd203;  #10 
a = 8'd107; b = 8'd204;  #10 
a = 8'd107; b = 8'd205;  #10 
a = 8'd107; b = 8'd206;  #10 
a = 8'd107; b = 8'd207;  #10 
a = 8'd107; b = 8'd208;  #10 
a = 8'd107; b = 8'd209;  #10 
a = 8'd107; b = 8'd210;  #10 
a = 8'd107; b = 8'd211;  #10 
a = 8'd107; b = 8'd212;  #10 
a = 8'd107; b = 8'd213;  #10 
a = 8'd107; b = 8'd214;  #10 
a = 8'd107; b = 8'd215;  #10 
a = 8'd107; b = 8'd216;  #10 
a = 8'd107; b = 8'd217;  #10 
a = 8'd107; b = 8'd218;  #10 
a = 8'd107; b = 8'd219;  #10 
a = 8'd107; b = 8'd220;  #10 
a = 8'd107; b = 8'd221;  #10 
a = 8'd107; b = 8'd222;  #10 
a = 8'd107; b = 8'd223;  #10 
a = 8'd107; b = 8'd224;  #10 
a = 8'd107; b = 8'd225;  #10 
a = 8'd107; b = 8'd226;  #10 
a = 8'd107; b = 8'd227;  #10 
a = 8'd107; b = 8'd228;  #10 
a = 8'd107; b = 8'd229;  #10 
a = 8'd107; b = 8'd230;  #10 
a = 8'd107; b = 8'd231;  #10 
a = 8'd107; b = 8'd232;  #10 
a = 8'd107; b = 8'd233;  #10 
a = 8'd107; b = 8'd234;  #10 
a = 8'd107; b = 8'd235;  #10 
a = 8'd107; b = 8'd236;  #10 
a = 8'd107; b = 8'd237;  #10 
a = 8'd107; b = 8'd238;  #10 
a = 8'd107; b = 8'd239;  #10 
a = 8'd107; b = 8'd240;  #10 
a = 8'd107; b = 8'd241;  #10 
a = 8'd107; b = 8'd242;  #10 
a = 8'd107; b = 8'd243;  #10 
a = 8'd107; b = 8'd244;  #10 
a = 8'd107; b = 8'd245;  #10 
a = 8'd107; b = 8'd246;  #10 
a = 8'd107; b = 8'd247;  #10 
a = 8'd107; b = 8'd248;  #10 
a = 8'd107; b = 8'd249;  #10 
a = 8'd107; b = 8'd250;  #10 
a = 8'd107; b = 8'd251;  #10 
a = 8'd107; b = 8'd252;  #10 
a = 8'd107; b = 8'd253;  #10 
a = 8'd107; b = 8'd254;  #10 
a = 8'd107; b = 8'd255;  #10 
a = 8'd108; b = 8'd0;  #10 
a = 8'd108; b = 8'd1;  #10 
a = 8'd108; b = 8'd2;  #10 
a = 8'd108; b = 8'd3;  #10 
a = 8'd108; b = 8'd4;  #10 
a = 8'd108; b = 8'd5;  #10 
a = 8'd108; b = 8'd6;  #10 
a = 8'd108; b = 8'd7;  #10 
a = 8'd108; b = 8'd8;  #10 
a = 8'd108; b = 8'd9;  #10 
a = 8'd108; b = 8'd10;  #10 
a = 8'd108; b = 8'd11;  #10 
a = 8'd108; b = 8'd12;  #10 
a = 8'd108; b = 8'd13;  #10 
a = 8'd108; b = 8'd14;  #10 
a = 8'd108; b = 8'd15;  #10 
a = 8'd108; b = 8'd16;  #10 
a = 8'd108; b = 8'd17;  #10 
a = 8'd108; b = 8'd18;  #10 
a = 8'd108; b = 8'd19;  #10 
a = 8'd108; b = 8'd20;  #10 
a = 8'd108; b = 8'd21;  #10 
a = 8'd108; b = 8'd22;  #10 
a = 8'd108; b = 8'd23;  #10 
a = 8'd108; b = 8'd24;  #10 
a = 8'd108; b = 8'd25;  #10 
a = 8'd108; b = 8'd26;  #10 
a = 8'd108; b = 8'd27;  #10 
a = 8'd108; b = 8'd28;  #10 
a = 8'd108; b = 8'd29;  #10 
a = 8'd108; b = 8'd30;  #10 
a = 8'd108; b = 8'd31;  #10 
a = 8'd108; b = 8'd32;  #10 
a = 8'd108; b = 8'd33;  #10 
a = 8'd108; b = 8'd34;  #10 
a = 8'd108; b = 8'd35;  #10 
a = 8'd108; b = 8'd36;  #10 
a = 8'd108; b = 8'd37;  #10 
a = 8'd108; b = 8'd38;  #10 
a = 8'd108; b = 8'd39;  #10 
a = 8'd108; b = 8'd40;  #10 
a = 8'd108; b = 8'd41;  #10 
a = 8'd108; b = 8'd42;  #10 
a = 8'd108; b = 8'd43;  #10 
a = 8'd108; b = 8'd44;  #10 
a = 8'd108; b = 8'd45;  #10 
a = 8'd108; b = 8'd46;  #10 
a = 8'd108; b = 8'd47;  #10 
a = 8'd108; b = 8'd48;  #10 
a = 8'd108; b = 8'd49;  #10 
a = 8'd108; b = 8'd50;  #10 
a = 8'd108; b = 8'd51;  #10 
a = 8'd108; b = 8'd52;  #10 
a = 8'd108; b = 8'd53;  #10 
a = 8'd108; b = 8'd54;  #10 
a = 8'd108; b = 8'd55;  #10 
a = 8'd108; b = 8'd56;  #10 
a = 8'd108; b = 8'd57;  #10 
a = 8'd108; b = 8'd58;  #10 
a = 8'd108; b = 8'd59;  #10 
a = 8'd108; b = 8'd60;  #10 
a = 8'd108; b = 8'd61;  #10 
a = 8'd108; b = 8'd62;  #10 
a = 8'd108; b = 8'd63;  #10 
a = 8'd108; b = 8'd64;  #10 
a = 8'd108; b = 8'd65;  #10 
a = 8'd108; b = 8'd66;  #10 
a = 8'd108; b = 8'd67;  #10 
a = 8'd108; b = 8'd68;  #10 
a = 8'd108; b = 8'd69;  #10 
a = 8'd108; b = 8'd70;  #10 
a = 8'd108; b = 8'd71;  #10 
a = 8'd108; b = 8'd72;  #10 
a = 8'd108; b = 8'd73;  #10 
a = 8'd108; b = 8'd74;  #10 
a = 8'd108; b = 8'd75;  #10 
a = 8'd108; b = 8'd76;  #10 
a = 8'd108; b = 8'd77;  #10 
a = 8'd108; b = 8'd78;  #10 
a = 8'd108; b = 8'd79;  #10 
a = 8'd108; b = 8'd80;  #10 
a = 8'd108; b = 8'd81;  #10 
a = 8'd108; b = 8'd82;  #10 
a = 8'd108; b = 8'd83;  #10 
a = 8'd108; b = 8'd84;  #10 
a = 8'd108; b = 8'd85;  #10 
a = 8'd108; b = 8'd86;  #10 
a = 8'd108; b = 8'd87;  #10 
a = 8'd108; b = 8'd88;  #10 
a = 8'd108; b = 8'd89;  #10 
a = 8'd108; b = 8'd90;  #10 
a = 8'd108; b = 8'd91;  #10 
a = 8'd108; b = 8'd92;  #10 
a = 8'd108; b = 8'd93;  #10 
a = 8'd108; b = 8'd94;  #10 
a = 8'd108; b = 8'd95;  #10 
a = 8'd108; b = 8'd96;  #10 
a = 8'd108; b = 8'd97;  #10 
a = 8'd108; b = 8'd98;  #10 
a = 8'd108; b = 8'd99;  #10 
a = 8'd108; b = 8'd100;  #10 
a = 8'd108; b = 8'd101;  #10 
a = 8'd108; b = 8'd102;  #10 
a = 8'd108; b = 8'd103;  #10 
a = 8'd108; b = 8'd104;  #10 
a = 8'd108; b = 8'd105;  #10 
a = 8'd108; b = 8'd106;  #10 
a = 8'd108; b = 8'd107;  #10 
a = 8'd108; b = 8'd108;  #10 
a = 8'd108; b = 8'd109;  #10 
a = 8'd108; b = 8'd110;  #10 
a = 8'd108; b = 8'd111;  #10 
a = 8'd108; b = 8'd112;  #10 
a = 8'd108; b = 8'd113;  #10 
a = 8'd108; b = 8'd114;  #10 
a = 8'd108; b = 8'd115;  #10 
a = 8'd108; b = 8'd116;  #10 
a = 8'd108; b = 8'd117;  #10 
a = 8'd108; b = 8'd118;  #10 
a = 8'd108; b = 8'd119;  #10 
a = 8'd108; b = 8'd120;  #10 
a = 8'd108; b = 8'd121;  #10 
a = 8'd108; b = 8'd122;  #10 
a = 8'd108; b = 8'd123;  #10 
a = 8'd108; b = 8'd124;  #10 
a = 8'd108; b = 8'd125;  #10 
a = 8'd108; b = 8'd126;  #10 
a = 8'd108; b = 8'd127;  #10 
a = 8'd108; b = 8'd128;  #10 
a = 8'd108; b = 8'd129;  #10 
a = 8'd108; b = 8'd130;  #10 
a = 8'd108; b = 8'd131;  #10 
a = 8'd108; b = 8'd132;  #10 
a = 8'd108; b = 8'd133;  #10 
a = 8'd108; b = 8'd134;  #10 
a = 8'd108; b = 8'd135;  #10 
a = 8'd108; b = 8'd136;  #10 
a = 8'd108; b = 8'd137;  #10 
a = 8'd108; b = 8'd138;  #10 
a = 8'd108; b = 8'd139;  #10 
a = 8'd108; b = 8'd140;  #10 
a = 8'd108; b = 8'd141;  #10 
a = 8'd108; b = 8'd142;  #10 
a = 8'd108; b = 8'd143;  #10 
a = 8'd108; b = 8'd144;  #10 
a = 8'd108; b = 8'd145;  #10 
a = 8'd108; b = 8'd146;  #10 
a = 8'd108; b = 8'd147;  #10 
a = 8'd108; b = 8'd148;  #10 
a = 8'd108; b = 8'd149;  #10 
a = 8'd108; b = 8'd150;  #10 
a = 8'd108; b = 8'd151;  #10 
a = 8'd108; b = 8'd152;  #10 
a = 8'd108; b = 8'd153;  #10 
a = 8'd108; b = 8'd154;  #10 
a = 8'd108; b = 8'd155;  #10 
a = 8'd108; b = 8'd156;  #10 
a = 8'd108; b = 8'd157;  #10 
a = 8'd108; b = 8'd158;  #10 
a = 8'd108; b = 8'd159;  #10 
a = 8'd108; b = 8'd160;  #10 
a = 8'd108; b = 8'd161;  #10 
a = 8'd108; b = 8'd162;  #10 
a = 8'd108; b = 8'd163;  #10 
a = 8'd108; b = 8'd164;  #10 
a = 8'd108; b = 8'd165;  #10 
a = 8'd108; b = 8'd166;  #10 
a = 8'd108; b = 8'd167;  #10 
a = 8'd108; b = 8'd168;  #10 
a = 8'd108; b = 8'd169;  #10 
a = 8'd108; b = 8'd170;  #10 
a = 8'd108; b = 8'd171;  #10 
a = 8'd108; b = 8'd172;  #10 
a = 8'd108; b = 8'd173;  #10 
a = 8'd108; b = 8'd174;  #10 
a = 8'd108; b = 8'd175;  #10 
a = 8'd108; b = 8'd176;  #10 
a = 8'd108; b = 8'd177;  #10 
a = 8'd108; b = 8'd178;  #10 
a = 8'd108; b = 8'd179;  #10 
a = 8'd108; b = 8'd180;  #10 
a = 8'd108; b = 8'd181;  #10 
a = 8'd108; b = 8'd182;  #10 
a = 8'd108; b = 8'd183;  #10 
a = 8'd108; b = 8'd184;  #10 
a = 8'd108; b = 8'd185;  #10 
a = 8'd108; b = 8'd186;  #10 
a = 8'd108; b = 8'd187;  #10 
a = 8'd108; b = 8'd188;  #10 
a = 8'd108; b = 8'd189;  #10 
a = 8'd108; b = 8'd190;  #10 
a = 8'd108; b = 8'd191;  #10 
a = 8'd108; b = 8'd192;  #10 
a = 8'd108; b = 8'd193;  #10 
a = 8'd108; b = 8'd194;  #10 
a = 8'd108; b = 8'd195;  #10 
a = 8'd108; b = 8'd196;  #10 
a = 8'd108; b = 8'd197;  #10 
a = 8'd108; b = 8'd198;  #10 
a = 8'd108; b = 8'd199;  #10 
a = 8'd108; b = 8'd200;  #10 
a = 8'd108; b = 8'd201;  #10 
a = 8'd108; b = 8'd202;  #10 
a = 8'd108; b = 8'd203;  #10 
a = 8'd108; b = 8'd204;  #10 
a = 8'd108; b = 8'd205;  #10 
a = 8'd108; b = 8'd206;  #10 
a = 8'd108; b = 8'd207;  #10 
a = 8'd108; b = 8'd208;  #10 
a = 8'd108; b = 8'd209;  #10 
a = 8'd108; b = 8'd210;  #10 
a = 8'd108; b = 8'd211;  #10 
a = 8'd108; b = 8'd212;  #10 
a = 8'd108; b = 8'd213;  #10 
a = 8'd108; b = 8'd214;  #10 
a = 8'd108; b = 8'd215;  #10 
a = 8'd108; b = 8'd216;  #10 
a = 8'd108; b = 8'd217;  #10 
a = 8'd108; b = 8'd218;  #10 
a = 8'd108; b = 8'd219;  #10 
a = 8'd108; b = 8'd220;  #10 
a = 8'd108; b = 8'd221;  #10 
a = 8'd108; b = 8'd222;  #10 
a = 8'd108; b = 8'd223;  #10 
a = 8'd108; b = 8'd224;  #10 
a = 8'd108; b = 8'd225;  #10 
a = 8'd108; b = 8'd226;  #10 
a = 8'd108; b = 8'd227;  #10 
a = 8'd108; b = 8'd228;  #10 
a = 8'd108; b = 8'd229;  #10 
a = 8'd108; b = 8'd230;  #10 
a = 8'd108; b = 8'd231;  #10 
a = 8'd108; b = 8'd232;  #10 
a = 8'd108; b = 8'd233;  #10 
a = 8'd108; b = 8'd234;  #10 
a = 8'd108; b = 8'd235;  #10 
a = 8'd108; b = 8'd236;  #10 
a = 8'd108; b = 8'd237;  #10 
a = 8'd108; b = 8'd238;  #10 
a = 8'd108; b = 8'd239;  #10 
a = 8'd108; b = 8'd240;  #10 
a = 8'd108; b = 8'd241;  #10 
a = 8'd108; b = 8'd242;  #10 
a = 8'd108; b = 8'd243;  #10 
a = 8'd108; b = 8'd244;  #10 
a = 8'd108; b = 8'd245;  #10 
a = 8'd108; b = 8'd246;  #10 
a = 8'd108; b = 8'd247;  #10 
a = 8'd108; b = 8'd248;  #10 
a = 8'd108; b = 8'd249;  #10 
a = 8'd108; b = 8'd250;  #10 
a = 8'd108; b = 8'd251;  #10 
a = 8'd108; b = 8'd252;  #10 
a = 8'd108; b = 8'd253;  #10 
a = 8'd108; b = 8'd254;  #10 
a = 8'd108; b = 8'd255;  #10 
a = 8'd109; b = 8'd0;  #10 
a = 8'd109; b = 8'd1;  #10 
a = 8'd109; b = 8'd2;  #10 
a = 8'd109; b = 8'd3;  #10 
a = 8'd109; b = 8'd4;  #10 
a = 8'd109; b = 8'd5;  #10 
a = 8'd109; b = 8'd6;  #10 
a = 8'd109; b = 8'd7;  #10 
a = 8'd109; b = 8'd8;  #10 
a = 8'd109; b = 8'd9;  #10 
a = 8'd109; b = 8'd10;  #10 
a = 8'd109; b = 8'd11;  #10 
a = 8'd109; b = 8'd12;  #10 
a = 8'd109; b = 8'd13;  #10 
a = 8'd109; b = 8'd14;  #10 
a = 8'd109; b = 8'd15;  #10 
a = 8'd109; b = 8'd16;  #10 
a = 8'd109; b = 8'd17;  #10 
a = 8'd109; b = 8'd18;  #10 
a = 8'd109; b = 8'd19;  #10 
a = 8'd109; b = 8'd20;  #10 
a = 8'd109; b = 8'd21;  #10 
a = 8'd109; b = 8'd22;  #10 
a = 8'd109; b = 8'd23;  #10 
a = 8'd109; b = 8'd24;  #10 
a = 8'd109; b = 8'd25;  #10 
a = 8'd109; b = 8'd26;  #10 
a = 8'd109; b = 8'd27;  #10 
a = 8'd109; b = 8'd28;  #10 
a = 8'd109; b = 8'd29;  #10 
a = 8'd109; b = 8'd30;  #10 
a = 8'd109; b = 8'd31;  #10 
a = 8'd109; b = 8'd32;  #10 
a = 8'd109; b = 8'd33;  #10 
a = 8'd109; b = 8'd34;  #10 
a = 8'd109; b = 8'd35;  #10 
a = 8'd109; b = 8'd36;  #10 
a = 8'd109; b = 8'd37;  #10 
a = 8'd109; b = 8'd38;  #10 
a = 8'd109; b = 8'd39;  #10 
a = 8'd109; b = 8'd40;  #10 
a = 8'd109; b = 8'd41;  #10 
a = 8'd109; b = 8'd42;  #10 
a = 8'd109; b = 8'd43;  #10 
a = 8'd109; b = 8'd44;  #10 
a = 8'd109; b = 8'd45;  #10 
a = 8'd109; b = 8'd46;  #10 
a = 8'd109; b = 8'd47;  #10 
a = 8'd109; b = 8'd48;  #10 
a = 8'd109; b = 8'd49;  #10 
a = 8'd109; b = 8'd50;  #10 
a = 8'd109; b = 8'd51;  #10 
a = 8'd109; b = 8'd52;  #10 
a = 8'd109; b = 8'd53;  #10 
a = 8'd109; b = 8'd54;  #10 
a = 8'd109; b = 8'd55;  #10 
a = 8'd109; b = 8'd56;  #10 
a = 8'd109; b = 8'd57;  #10 
a = 8'd109; b = 8'd58;  #10 
a = 8'd109; b = 8'd59;  #10 
a = 8'd109; b = 8'd60;  #10 
a = 8'd109; b = 8'd61;  #10 
a = 8'd109; b = 8'd62;  #10 
a = 8'd109; b = 8'd63;  #10 
a = 8'd109; b = 8'd64;  #10 
a = 8'd109; b = 8'd65;  #10 
a = 8'd109; b = 8'd66;  #10 
a = 8'd109; b = 8'd67;  #10 
a = 8'd109; b = 8'd68;  #10 
a = 8'd109; b = 8'd69;  #10 
a = 8'd109; b = 8'd70;  #10 
a = 8'd109; b = 8'd71;  #10 
a = 8'd109; b = 8'd72;  #10 
a = 8'd109; b = 8'd73;  #10 
a = 8'd109; b = 8'd74;  #10 
a = 8'd109; b = 8'd75;  #10 
a = 8'd109; b = 8'd76;  #10 
a = 8'd109; b = 8'd77;  #10 
a = 8'd109; b = 8'd78;  #10 
a = 8'd109; b = 8'd79;  #10 
a = 8'd109; b = 8'd80;  #10 
a = 8'd109; b = 8'd81;  #10 
a = 8'd109; b = 8'd82;  #10 
a = 8'd109; b = 8'd83;  #10 
a = 8'd109; b = 8'd84;  #10 
a = 8'd109; b = 8'd85;  #10 
a = 8'd109; b = 8'd86;  #10 
a = 8'd109; b = 8'd87;  #10 
a = 8'd109; b = 8'd88;  #10 
a = 8'd109; b = 8'd89;  #10 
a = 8'd109; b = 8'd90;  #10 
a = 8'd109; b = 8'd91;  #10 
a = 8'd109; b = 8'd92;  #10 
a = 8'd109; b = 8'd93;  #10 
a = 8'd109; b = 8'd94;  #10 
a = 8'd109; b = 8'd95;  #10 
a = 8'd109; b = 8'd96;  #10 
a = 8'd109; b = 8'd97;  #10 
a = 8'd109; b = 8'd98;  #10 
a = 8'd109; b = 8'd99;  #10 
a = 8'd109; b = 8'd100;  #10 
a = 8'd109; b = 8'd101;  #10 
a = 8'd109; b = 8'd102;  #10 
a = 8'd109; b = 8'd103;  #10 
a = 8'd109; b = 8'd104;  #10 
a = 8'd109; b = 8'd105;  #10 
a = 8'd109; b = 8'd106;  #10 
a = 8'd109; b = 8'd107;  #10 
a = 8'd109; b = 8'd108;  #10 
a = 8'd109; b = 8'd109;  #10 
a = 8'd109; b = 8'd110;  #10 
a = 8'd109; b = 8'd111;  #10 
a = 8'd109; b = 8'd112;  #10 
a = 8'd109; b = 8'd113;  #10 
a = 8'd109; b = 8'd114;  #10 
a = 8'd109; b = 8'd115;  #10 
a = 8'd109; b = 8'd116;  #10 
a = 8'd109; b = 8'd117;  #10 
a = 8'd109; b = 8'd118;  #10 
a = 8'd109; b = 8'd119;  #10 
a = 8'd109; b = 8'd120;  #10 
a = 8'd109; b = 8'd121;  #10 
a = 8'd109; b = 8'd122;  #10 
a = 8'd109; b = 8'd123;  #10 
a = 8'd109; b = 8'd124;  #10 
a = 8'd109; b = 8'd125;  #10 
a = 8'd109; b = 8'd126;  #10 
a = 8'd109; b = 8'd127;  #10 
a = 8'd109; b = 8'd128;  #10 
a = 8'd109; b = 8'd129;  #10 
a = 8'd109; b = 8'd130;  #10 
a = 8'd109; b = 8'd131;  #10 
a = 8'd109; b = 8'd132;  #10 
a = 8'd109; b = 8'd133;  #10 
a = 8'd109; b = 8'd134;  #10 
a = 8'd109; b = 8'd135;  #10 
a = 8'd109; b = 8'd136;  #10 
a = 8'd109; b = 8'd137;  #10 
a = 8'd109; b = 8'd138;  #10 
a = 8'd109; b = 8'd139;  #10 
a = 8'd109; b = 8'd140;  #10 
a = 8'd109; b = 8'd141;  #10 
a = 8'd109; b = 8'd142;  #10 
a = 8'd109; b = 8'd143;  #10 
a = 8'd109; b = 8'd144;  #10 
a = 8'd109; b = 8'd145;  #10 
a = 8'd109; b = 8'd146;  #10 
a = 8'd109; b = 8'd147;  #10 
a = 8'd109; b = 8'd148;  #10 
a = 8'd109; b = 8'd149;  #10 
a = 8'd109; b = 8'd150;  #10 
a = 8'd109; b = 8'd151;  #10 
a = 8'd109; b = 8'd152;  #10 
a = 8'd109; b = 8'd153;  #10 
a = 8'd109; b = 8'd154;  #10 
a = 8'd109; b = 8'd155;  #10 
a = 8'd109; b = 8'd156;  #10 
a = 8'd109; b = 8'd157;  #10 
a = 8'd109; b = 8'd158;  #10 
a = 8'd109; b = 8'd159;  #10 
a = 8'd109; b = 8'd160;  #10 
a = 8'd109; b = 8'd161;  #10 
a = 8'd109; b = 8'd162;  #10 
a = 8'd109; b = 8'd163;  #10 
a = 8'd109; b = 8'd164;  #10 
a = 8'd109; b = 8'd165;  #10 
a = 8'd109; b = 8'd166;  #10 
a = 8'd109; b = 8'd167;  #10 
a = 8'd109; b = 8'd168;  #10 
a = 8'd109; b = 8'd169;  #10 
a = 8'd109; b = 8'd170;  #10 
a = 8'd109; b = 8'd171;  #10 
a = 8'd109; b = 8'd172;  #10 
a = 8'd109; b = 8'd173;  #10 
a = 8'd109; b = 8'd174;  #10 
a = 8'd109; b = 8'd175;  #10 
a = 8'd109; b = 8'd176;  #10 
a = 8'd109; b = 8'd177;  #10 
a = 8'd109; b = 8'd178;  #10 
a = 8'd109; b = 8'd179;  #10 
a = 8'd109; b = 8'd180;  #10 
a = 8'd109; b = 8'd181;  #10 
a = 8'd109; b = 8'd182;  #10 
a = 8'd109; b = 8'd183;  #10 
a = 8'd109; b = 8'd184;  #10 
a = 8'd109; b = 8'd185;  #10 
a = 8'd109; b = 8'd186;  #10 
a = 8'd109; b = 8'd187;  #10 
a = 8'd109; b = 8'd188;  #10 
a = 8'd109; b = 8'd189;  #10 
a = 8'd109; b = 8'd190;  #10 
a = 8'd109; b = 8'd191;  #10 
a = 8'd109; b = 8'd192;  #10 
a = 8'd109; b = 8'd193;  #10 
a = 8'd109; b = 8'd194;  #10 
a = 8'd109; b = 8'd195;  #10 
a = 8'd109; b = 8'd196;  #10 
a = 8'd109; b = 8'd197;  #10 
a = 8'd109; b = 8'd198;  #10 
a = 8'd109; b = 8'd199;  #10 
a = 8'd109; b = 8'd200;  #10 
a = 8'd109; b = 8'd201;  #10 
a = 8'd109; b = 8'd202;  #10 
a = 8'd109; b = 8'd203;  #10 
a = 8'd109; b = 8'd204;  #10 
a = 8'd109; b = 8'd205;  #10 
a = 8'd109; b = 8'd206;  #10 
a = 8'd109; b = 8'd207;  #10 
a = 8'd109; b = 8'd208;  #10 
a = 8'd109; b = 8'd209;  #10 
a = 8'd109; b = 8'd210;  #10 
a = 8'd109; b = 8'd211;  #10 
a = 8'd109; b = 8'd212;  #10 
a = 8'd109; b = 8'd213;  #10 
a = 8'd109; b = 8'd214;  #10 
a = 8'd109; b = 8'd215;  #10 
a = 8'd109; b = 8'd216;  #10 
a = 8'd109; b = 8'd217;  #10 
a = 8'd109; b = 8'd218;  #10 
a = 8'd109; b = 8'd219;  #10 
a = 8'd109; b = 8'd220;  #10 
a = 8'd109; b = 8'd221;  #10 
a = 8'd109; b = 8'd222;  #10 
a = 8'd109; b = 8'd223;  #10 
a = 8'd109; b = 8'd224;  #10 
a = 8'd109; b = 8'd225;  #10 
a = 8'd109; b = 8'd226;  #10 
a = 8'd109; b = 8'd227;  #10 
a = 8'd109; b = 8'd228;  #10 
a = 8'd109; b = 8'd229;  #10 
a = 8'd109; b = 8'd230;  #10 
a = 8'd109; b = 8'd231;  #10 
a = 8'd109; b = 8'd232;  #10 
a = 8'd109; b = 8'd233;  #10 
a = 8'd109; b = 8'd234;  #10 
a = 8'd109; b = 8'd235;  #10 
a = 8'd109; b = 8'd236;  #10 
a = 8'd109; b = 8'd237;  #10 
a = 8'd109; b = 8'd238;  #10 
a = 8'd109; b = 8'd239;  #10 
a = 8'd109; b = 8'd240;  #10 
a = 8'd109; b = 8'd241;  #10 
a = 8'd109; b = 8'd242;  #10 
a = 8'd109; b = 8'd243;  #10 
a = 8'd109; b = 8'd244;  #10 
a = 8'd109; b = 8'd245;  #10 
a = 8'd109; b = 8'd246;  #10 
a = 8'd109; b = 8'd247;  #10 
a = 8'd109; b = 8'd248;  #10 
a = 8'd109; b = 8'd249;  #10 
a = 8'd109; b = 8'd250;  #10 
a = 8'd109; b = 8'd251;  #10 
a = 8'd109; b = 8'd252;  #10 
a = 8'd109; b = 8'd253;  #10 
a = 8'd109; b = 8'd254;  #10 
a = 8'd109; b = 8'd255;  #10 
a = 8'd110; b = 8'd0;  #10 
a = 8'd110; b = 8'd1;  #10 
a = 8'd110; b = 8'd2;  #10 
a = 8'd110; b = 8'd3;  #10 
a = 8'd110; b = 8'd4;  #10 
a = 8'd110; b = 8'd5;  #10 
a = 8'd110; b = 8'd6;  #10 
a = 8'd110; b = 8'd7;  #10 
a = 8'd110; b = 8'd8;  #10 
a = 8'd110; b = 8'd9;  #10 
a = 8'd110; b = 8'd10;  #10 
a = 8'd110; b = 8'd11;  #10 
a = 8'd110; b = 8'd12;  #10 
a = 8'd110; b = 8'd13;  #10 
a = 8'd110; b = 8'd14;  #10 
a = 8'd110; b = 8'd15;  #10 
a = 8'd110; b = 8'd16;  #10 
a = 8'd110; b = 8'd17;  #10 
a = 8'd110; b = 8'd18;  #10 
a = 8'd110; b = 8'd19;  #10 
a = 8'd110; b = 8'd20;  #10 
a = 8'd110; b = 8'd21;  #10 
a = 8'd110; b = 8'd22;  #10 
a = 8'd110; b = 8'd23;  #10 
a = 8'd110; b = 8'd24;  #10 
a = 8'd110; b = 8'd25;  #10 
a = 8'd110; b = 8'd26;  #10 
a = 8'd110; b = 8'd27;  #10 
a = 8'd110; b = 8'd28;  #10 
a = 8'd110; b = 8'd29;  #10 
a = 8'd110; b = 8'd30;  #10 
a = 8'd110; b = 8'd31;  #10 
a = 8'd110; b = 8'd32;  #10 
a = 8'd110; b = 8'd33;  #10 
a = 8'd110; b = 8'd34;  #10 
a = 8'd110; b = 8'd35;  #10 
a = 8'd110; b = 8'd36;  #10 
a = 8'd110; b = 8'd37;  #10 
a = 8'd110; b = 8'd38;  #10 
a = 8'd110; b = 8'd39;  #10 
a = 8'd110; b = 8'd40;  #10 
a = 8'd110; b = 8'd41;  #10 
a = 8'd110; b = 8'd42;  #10 
a = 8'd110; b = 8'd43;  #10 
a = 8'd110; b = 8'd44;  #10 
a = 8'd110; b = 8'd45;  #10 
a = 8'd110; b = 8'd46;  #10 
a = 8'd110; b = 8'd47;  #10 
a = 8'd110; b = 8'd48;  #10 
a = 8'd110; b = 8'd49;  #10 
a = 8'd110; b = 8'd50;  #10 
a = 8'd110; b = 8'd51;  #10 
a = 8'd110; b = 8'd52;  #10 
a = 8'd110; b = 8'd53;  #10 
a = 8'd110; b = 8'd54;  #10 
a = 8'd110; b = 8'd55;  #10 
a = 8'd110; b = 8'd56;  #10 
a = 8'd110; b = 8'd57;  #10 
a = 8'd110; b = 8'd58;  #10 
a = 8'd110; b = 8'd59;  #10 
a = 8'd110; b = 8'd60;  #10 
a = 8'd110; b = 8'd61;  #10 
a = 8'd110; b = 8'd62;  #10 
a = 8'd110; b = 8'd63;  #10 
a = 8'd110; b = 8'd64;  #10 
a = 8'd110; b = 8'd65;  #10 
a = 8'd110; b = 8'd66;  #10 
a = 8'd110; b = 8'd67;  #10 
a = 8'd110; b = 8'd68;  #10 
a = 8'd110; b = 8'd69;  #10 
a = 8'd110; b = 8'd70;  #10 
a = 8'd110; b = 8'd71;  #10 
a = 8'd110; b = 8'd72;  #10 
a = 8'd110; b = 8'd73;  #10 
a = 8'd110; b = 8'd74;  #10 
a = 8'd110; b = 8'd75;  #10 
a = 8'd110; b = 8'd76;  #10 
a = 8'd110; b = 8'd77;  #10 
a = 8'd110; b = 8'd78;  #10 
a = 8'd110; b = 8'd79;  #10 
a = 8'd110; b = 8'd80;  #10 
a = 8'd110; b = 8'd81;  #10 
a = 8'd110; b = 8'd82;  #10 
a = 8'd110; b = 8'd83;  #10 
a = 8'd110; b = 8'd84;  #10 
a = 8'd110; b = 8'd85;  #10 
a = 8'd110; b = 8'd86;  #10 
a = 8'd110; b = 8'd87;  #10 
a = 8'd110; b = 8'd88;  #10 
a = 8'd110; b = 8'd89;  #10 
a = 8'd110; b = 8'd90;  #10 
a = 8'd110; b = 8'd91;  #10 
a = 8'd110; b = 8'd92;  #10 
a = 8'd110; b = 8'd93;  #10 
a = 8'd110; b = 8'd94;  #10 
a = 8'd110; b = 8'd95;  #10 
a = 8'd110; b = 8'd96;  #10 
a = 8'd110; b = 8'd97;  #10 
a = 8'd110; b = 8'd98;  #10 
a = 8'd110; b = 8'd99;  #10 
a = 8'd110; b = 8'd100;  #10 
a = 8'd110; b = 8'd101;  #10 
a = 8'd110; b = 8'd102;  #10 
a = 8'd110; b = 8'd103;  #10 
a = 8'd110; b = 8'd104;  #10 
a = 8'd110; b = 8'd105;  #10 
a = 8'd110; b = 8'd106;  #10 
a = 8'd110; b = 8'd107;  #10 
a = 8'd110; b = 8'd108;  #10 
a = 8'd110; b = 8'd109;  #10 
a = 8'd110; b = 8'd110;  #10 
a = 8'd110; b = 8'd111;  #10 
a = 8'd110; b = 8'd112;  #10 
a = 8'd110; b = 8'd113;  #10 
a = 8'd110; b = 8'd114;  #10 
a = 8'd110; b = 8'd115;  #10 
a = 8'd110; b = 8'd116;  #10 
a = 8'd110; b = 8'd117;  #10 
a = 8'd110; b = 8'd118;  #10 
a = 8'd110; b = 8'd119;  #10 
a = 8'd110; b = 8'd120;  #10 
a = 8'd110; b = 8'd121;  #10 
a = 8'd110; b = 8'd122;  #10 
a = 8'd110; b = 8'd123;  #10 
a = 8'd110; b = 8'd124;  #10 
a = 8'd110; b = 8'd125;  #10 
a = 8'd110; b = 8'd126;  #10 
a = 8'd110; b = 8'd127;  #10 
a = 8'd110; b = 8'd128;  #10 
a = 8'd110; b = 8'd129;  #10 
a = 8'd110; b = 8'd130;  #10 
a = 8'd110; b = 8'd131;  #10 
a = 8'd110; b = 8'd132;  #10 
a = 8'd110; b = 8'd133;  #10 
a = 8'd110; b = 8'd134;  #10 
a = 8'd110; b = 8'd135;  #10 
a = 8'd110; b = 8'd136;  #10 
a = 8'd110; b = 8'd137;  #10 
a = 8'd110; b = 8'd138;  #10 
a = 8'd110; b = 8'd139;  #10 
a = 8'd110; b = 8'd140;  #10 
a = 8'd110; b = 8'd141;  #10 
a = 8'd110; b = 8'd142;  #10 
a = 8'd110; b = 8'd143;  #10 
a = 8'd110; b = 8'd144;  #10 
a = 8'd110; b = 8'd145;  #10 
a = 8'd110; b = 8'd146;  #10 
a = 8'd110; b = 8'd147;  #10 
a = 8'd110; b = 8'd148;  #10 
a = 8'd110; b = 8'd149;  #10 
a = 8'd110; b = 8'd150;  #10 
a = 8'd110; b = 8'd151;  #10 
a = 8'd110; b = 8'd152;  #10 
a = 8'd110; b = 8'd153;  #10 
a = 8'd110; b = 8'd154;  #10 
a = 8'd110; b = 8'd155;  #10 
a = 8'd110; b = 8'd156;  #10 
a = 8'd110; b = 8'd157;  #10 
a = 8'd110; b = 8'd158;  #10 
a = 8'd110; b = 8'd159;  #10 
a = 8'd110; b = 8'd160;  #10 
a = 8'd110; b = 8'd161;  #10 
a = 8'd110; b = 8'd162;  #10 
a = 8'd110; b = 8'd163;  #10 
a = 8'd110; b = 8'd164;  #10 
a = 8'd110; b = 8'd165;  #10 
a = 8'd110; b = 8'd166;  #10 
a = 8'd110; b = 8'd167;  #10 
a = 8'd110; b = 8'd168;  #10 
a = 8'd110; b = 8'd169;  #10 
a = 8'd110; b = 8'd170;  #10 
a = 8'd110; b = 8'd171;  #10 
a = 8'd110; b = 8'd172;  #10 
a = 8'd110; b = 8'd173;  #10 
a = 8'd110; b = 8'd174;  #10 
a = 8'd110; b = 8'd175;  #10 
a = 8'd110; b = 8'd176;  #10 
a = 8'd110; b = 8'd177;  #10 
a = 8'd110; b = 8'd178;  #10 
a = 8'd110; b = 8'd179;  #10 
a = 8'd110; b = 8'd180;  #10 
a = 8'd110; b = 8'd181;  #10 
a = 8'd110; b = 8'd182;  #10 
a = 8'd110; b = 8'd183;  #10 
a = 8'd110; b = 8'd184;  #10 
a = 8'd110; b = 8'd185;  #10 
a = 8'd110; b = 8'd186;  #10 
a = 8'd110; b = 8'd187;  #10 
a = 8'd110; b = 8'd188;  #10 
a = 8'd110; b = 8'd189;  #10 
a = 8'd110; b = 8'd190;  #10 
a = 8'd110; b = 8'd191;  #10 
a = 8'd110; b = 8'd192;  #10 
a = 8'd110; b = 8'd193;  #10 
a = 8'd110; b = 8'd194;  #10 
a = 8'd110; b = 8'd195;  #10 
a = 8'd110; b = 8'd196;  #10 
a = 8'd110; b = 8'd197;  #10 
a = 8'd110; b = 8'd198;  #10 
a = 8'd110; b = 8'd199;  #10 
a = 8'd110; b = 8'd200;  #10 
a = 8'd110; b = 8'd201;  #10 
a = 8'd110; b = 8'd202;  #10 
a = 8'd110; b = 8'd203;  #10 
a = 8'd110; b = 8'd204;  #10 
a = 8'd110; b = 8'd205;  #10 
a = 8'd110; b = 8'd206;  #10 
a = 8'd110; b = 8'd207;  #10 
a = 8'd110; b = 8'd208;  #10 
a = 8'd110; b = 8'd209;  #10 
a = 8'd110; b = 8'd210;  #10 
a = 8'd110; b = 8'd211;  #10 
a = 8'd110; b = 8'd212;  #10 
a = 8'd110; b = 8'd213;  #10 
a = 8'd110; b = 8'd214;  #10 
a = 8'd110; b = 8'd215;  #10 
a = 8'd110; b = 8'd216;  #10 
a = 8'd110; b = 8'd217;  #10 
a = 8'd110; b = 8'd218;  #10 
a = 8'd110; b = 8'd219;  #10 
a = 8'd110; b = 8'd220;  #10 
a = 8'd110; b = 8'd221;  #10 
a = 8'd110; b = 8'd222;  #10 
a = 8'd110; b = 8'd223;  #10 
a = 8'd110; b = 8'd224;  #10 
a = 8'd110; b = 8'd225;  #10 
a = 8'd110; b = 8'd226;  #10 
a = 8'd110; b = 8'd227;  #10 
a = 8'd110; b = 8'd228;  #10 
a = 8'd110; b = 8'd229;  #10 
a = 8'd110; b = 8'd230;  #10 
a = 8'd110; b = 8'd231;  #10 
a = 8'd110; b = 8'd232;  #10 
a = 8'd110; b = 8'd233;  #10 
a = 8'd110; b = 8'd234;  #10 
a = 8'd110; b = 8'd235;  #10 
a = 8'd110; b = 8'd236;  #10 
a = 8'd110; b = 8'd237;  #10 
a = 8'd110; b = 8'd238;  #10 
a = 8'd110; b = 8'd239;  #10 
a = 8'd110; b = 8'd240;  #10 
a = 8'd110; b = 8'd241;  #10 
a = 8'd110; b = 8'd242;  #10 
a = 8'd110; b = 8'd243;  #10 
a = 8'd110; b = 8'd244;  #10 
a = 8'd110; b = 8'd245;  #10 
a = 8'd110; b = 8'd246;  #10 
a = 8'd110; b = 8'd247;  #10 
a = 8'd110; b = 8'd248;  #10 
a = 8'd110; b = 8'd249;  #10 
a = 8'd110; b = 8'd250;  #10 
a = 8'd110; b = 8'd251;  #10 
a = 8'd110; b = 8'd252;  #10 
a = 8'd110; b = 8'd253;  #10 
a = 8'd110; b = 8'd254;  #10 
a = 8'd110; b = 8'd255;  #10 
a = 8'd111; b = 8'd0;  #10 
a = 8'd111; b = 8'd1;  #10 
a = 8'd111; b = 8'd2;  #10 
a = 8'd111; b = 8'd3;  #10 
a = 8'd111; b = 8'd4;  #10 
a = 8'd111; b = 8'd5;  #10 
a = 8'd111; b = 8'd6;  #10 
a = 8'd111; b = 8'd7;  #10 
a = 8'd111; b = 8'd8;  #10 
a = 8'd111; b = 8'd9;  #10 
a = 8'd111; b = 8'd10;  #10 
a = 8'd111; b = 8'd11;  #10 
a = 8'd111; b = 8'd12;  #10 
a = 8'd111; b = 8'd13;  #10 
a = 8'd111; b = 8'd14;  #10 
a = 8'd111; b = 8'd15;  #10 
a = 8'd111; b = 8'd16;  #10 
a = 8'd111; b = 8'd17;  #10 
a = 8'd111; b = 8'd18;  #10 
a = 8'd111; b = 8'd19;  #10 
a = 8'd111; b = 8'd20;  #10 
a = 8'd111; b = 8'd21;  #10 
a = 8'd111; b = 8'd22;  #10 
a = 8'd111; b = 8'd23;  #10 
a = 8'd111; b = 8'd24;  #10 
a = 8'd111; b = 8'd25;  #10 
a = 8'd111; b = 8'd26;  #10 
a = 8'd111; b = 8'd27;  #10 
a = 8'd111; b = 8'd28;  #10 
a = 8'd111; b = 8'd29;  #10 
a = 8'd111; b = 8'd30;  #10 
a = 8'd111; b = 8'd31;  #10 
a = 8'd111; b = 8'd32;  #10 
a = 8'd111; b = 8'd33;  #10 
a = 8'd111; b = 8'd34;  #10 
a = 8'd111; b = 8'd35;  #10 
a = 8'd111; b = 8'd36;  #10 
a = 8'd111; b = 8'd37;  #10 
a = 8'd111; b = 8'd38;  #10 
a = 8'd111; b = 8'd39;  #10 
a = 8'd111; b = 8'd40;  #10 
a = 8'd111; b = 8'd41;  #10 
a = 8'd111; b = 8'd42;  #10 
a = 8'd111; b = 8'd43;  #10 
a = 8'd111; b = 8'd44;  #10 
a = 8'd111; b = 8'd45;  #10 
a = 8'd111; b = 8'd46;  #10 
a = 8'd111; b = 8'd47;  #10 
a = 8'd111; b = 8'd48;  #10 
a = 8'd111; b = 8'd49;  #10 
a = 8'd111; b = 8'd50;  #10 
a = 8'd111; b = 8'd51;  #10 
a = 8'd111; b = 8'd52;  #10 
a = 8'd111; b = 8'd53;  #10 
a = 8'd111; b = 8'd54;  #10 
a = 8'd111; b = 8'd55;  #10 
a = 8'd111; b = 8'd56;  #10 
a = 8'd111; b = 8'd57;  #10 
a = 8'd111; b = 8'd58;  #10 
a = 8'd111; b = 8'd59;  #10 
a = 8'd111; b = 8'd60;  #10 
a = 8'd111; b = 8'd61;  #10 
a = 8'd111; b = 8'd62;  #10 
a = 8'd111; b = 8'd63;  #10 
a = 8'd111; b = 8'd64;  #10 
a = 8'd111; b = 8'd65;  #10 
a = 8'd111; b = 8'd66;  #10 
a = 8'd111; b = 8'd67;  #10 
a = 8'd111; b = 8'd68;  #10 
a = 8'd111; b = 8'd69;  #10 
a = 8'd111; b = 8'd70;  #10 
a = 8'd111; b = 8'd71;  #10 
a = 8'd111; b = 8'd72;  #10 
a = 8'd111; b = 8'd73;  #10 
a = 8'd111; b = 8'd74;  #10 
a = 8'd111; b = 8'd75;  #10 
a = 8'd111; b = 8'd76;  #10 
a = 8'd111; b = 8'd77;  #10 
a = 8'd111; b = 8'd78;  #10 
a = 8'd111; b = 8'd79;  #10 
a = 8'd111; b = 8'd80;  #10 
a = 8'd111; b = 8'd81;  #10 
a = 8'd111; b = 8'd82;  #10 
a = 8'd111; b = 8'd83;  #10 
a = 8'd111; b = 8'd84;  #10 
a = 8'd111; b = 8'd85;  #10 
a = 8'd111; b = 8'd86;  #10 
a = 8'd111; b = 8'd87;  #10 
a = 8'd111; b = 8'd88;  #10 
a = 8'd111; b = 8'd89;  #10 
a = 8'd111; b = 8'd90;  #10 
a = 8'd111; b = 8'd91;  #10 
a = 8'd111; b = 8'd92;  #10 
a = 8'd111; b = 8'd93;  #10 
a = 8'd111; b = 8'd94;  #10 
a = 8'd111; b = 8'd95;  #10 
a = 8'd111; b = 8'd96;  #10 
a = 8'd111; b = 8'd97;  #10 
a = 8'd111; b = 8'd98;  #10 
a = 8'd111; b = 8'd99;  #10 
a = 8'd111; b = 8'd100;  #10 
a = 8'd111; b = 8'd101;  #10 
a = 8'd111; b = 8'd102;  #10 
a = 8'd111; b = 8'd103;  #10 
a = 8'd111; b = 8'd104;  #10 
a = 8'd111; b = 8'd105;  #10 
a = 8'd111; b = 8'd106;  #10 
a = 8'd111; b = 8'd107;  #10 
a = 8'd111; b = 8'd108;  #10 
a = 8'd111; b = 8'd109;  #10 
a = 8'd111; b = 8'd110;  #10 
a = 8'd111; b = 8'd111;  #10 
a = 8'd111; b = 8'd112;  #10 
a = 8'd111; b = 8'd113;  #10 
a = 8'd111; b = 8'd114;  #10 
a = 8'd111; b = 8'd115;  #10 
a = 8'd111; b = 8'd116;  #10 
a = 8'd111; b = 8'd117;  #10 
a = 8'd111; b = 8'd118;  #10 
a = 8'd111; b = 8'd119;  #10 
a = 8'd111; b = 8'd120;  #10 
a = 8'd111; b = 8'd121;  #10 
a = 8'd111; b = 8'd122;  #10 
a = 8'd111; b = 8'd123;  #10 
a = 8'd111; b = 8'd124;  #10 
a = 8'd111; b = 8'd125;  #10 
a = 8'd111; b = 8'd126;  #10 
a = 8'd111; b = 8'd127;  #10 
a = 8'd111; b = 8'd128;  #10 
a = 8'd111; b = 8'd129;  #10 
a = 8'd111; b = 8'd130;  #10 
a = 8'd111; b = 8'd131;  #10 
a = 8'd111; b = 8'd132;  #10 
a = 8'd111; b = 8'd133;  #10 
a = 8'd111; b = 8'd134;  #10 
a = 8'd111; b = 8'd135;  #10 
a = 8'd111; b = 8'd136;  #10 
a = 8'd111; b = 8'd137;  #10 
a = 8'd111; b = 8'd138;  #10 
a = 8'd111; b = 8'd139;  #10 
a = 8'd111; b = 8'd140;  #10 
a = 8'd111; b = 8'd141;  #10 
a = 8'd111; b = 8'd142;  #10 
a = 8'd111; b = 8'd143;  #10 
a = 8'd111; b = 8'd144;  #10 
a = 8'd111; b = 8'd145;  #10 
a = 8'd111; b = 8'd146;  #10 
a = 8'd111; b = 8'd147;  #10 
a = 8'd111; b = 8'd148;  #10 
a = 8'd111; b = 8'd149;  #10 
a = 8'd111; b = 8'd150;  #10 
a = 8'd111; b = 8'd151;  #10 
a = 8'd111; b = 8'd152;  #10 
a = 8'd111; b = 8'd153;  #10 
a = 8'd111; b = 8'd154;  #10 
a = 8'd111; b = 8'd155;  #10 
a = 8'd111; b = 8'd156;  #10 
a = 8'd111; b = 8'd157;  #10 
a = 8'd111; b = 8'd158;  #10 
a = 8'd111; b = 8'd159;  #10 
a = 8'd111; b = 8'd160;  #10 
a = 8'd111; b = 8'd161;  #10 
a = 8'd111; b = 8'd162;  #10 
a = 8'd111; b = 8'd163;  #10 
a = 8'd111; b = 8'd164;  #10 
a = 8'd111; b = 8'd165;  #10 
a = 8'd111; b = 8'd166;  #10 
a = 8'd111; b = 8'd167;  #10 
a = 8'd111; b = 8'd168;  #10 
a = 8'd111; b = 8'd169;  #10 
a = 8'd111; b = 8'd170;  #10 
a = 8'd111; b = 8'd171;  #10 
a = 8'd111; b = 8'd172;  #10 
a = 8'd111; b = 8'd173;  #10 
a = 8'd111; b = 8'd174;  #10 
a = 8'd111; b = 8'd175;  #10 
a = 8'd111; b = 8'd176;  #10 
a = 8'd111; b = 8'd177;  #10 
a = 8'd111; b = 8'd178;  #10 
a = 8'd111; b = 8'd179;  #10 
a = 8'd111; b = 8'd180;  #10 
a = 8'd111; b = 8'd181;  #10 
a = 8'd111; b = 8'd182;  #10 
a = 8'd111; b = 8'd183;  #10 
a = 8'd111; b = 8'd184;  #10 
a = 8'd111; b = 8'd185;  #10 
a = 8'd111; b = 8'd186;  #10 
a = 8'd111; b = 8'd187;  #10 
a = 8'd111; b = 8'd188;  #10 
a = 8'd111; b = 8'd189;  #10 
a = 8'd111; b = 8'd190;  #10 
a = 8'd111; b = 8'd191;  #10 
a = 8'd111; b = 8'd192;  #10 
a = 8'd111; b = 8'd193;  #10 
a = 8'd111; b = 8'd194;  #10 
a = 8'd111; b = 8'd195;  #10 
a = 8'd111; b = 8'd196;  #10 
a = 8'd111; b = 8'd197;  #10 
a = 8'd111; b = 8'd198;  #10 
a = 8'd111; b = 8'd199;  #10 
a = 8'd111; b = 8'd200;  #10 
a = 8'd111; b = 8'd201;  #10 
a = 8'd111; b = 8'd202;  #10 
a = 8'd111; b = 8'd203;  #10 
a = 8'd111; b = 8'd204;  #10 
a = 8'd111; b = 8'd205;  #10 
a = 8'd111; b = 8'd206;  #10 
a = 8'd111; b = 8'd207;  #10 
a = 8'd111; b = 8'd208;  #10 
a = 8'd111; b = 8'd209;  #10 
a = 8'd111; b = 8'd210;  #10 
a = 8'd111; b = 8'd211;  #10 
a = 8'd111; b = 8'd212;  #10 
a = 8'd111; b = 8'd213;  #10 
a = 8'd111; b = 8'd214;  #10 
a = 8'd111; b = 8'd215;  #10 
a = 8'd111; b = 8'd216;  #10 
a = 8'd111; b = 8'd217;  #10 
a = 8'd111; b = 8'd218;  #10 
a = 8'd111; b = 8'd219;  #10 
a = 8'd111; b = 8'd220;  #10 
a = 8'd111; b = 8'd221;  #10 
a = 8'd111; b = 8'd222;  #10 
a = 8'd111; b = 8'd223;  #10 
a = 8'd111; b = 8'd224;  #10 
a = 8'd111; b = 8'd225;  #10 
a = 8'd111; b = 8'd226;  #10 
a = 8'd111; b = 8'd227;  #10 
a = 8'd111; b = 8'd228;  #10 
a = 8'd111; b = 8'd229;  #10 
a = 8'd111; b = 8'd230;  #10 
a = 8'd111; b = 8'd231;  #10 
a = 8'd111; b = 8'd232;  #10 
a = 8'd111; b = 8'd233;  #10 
a = 8'd111; b = 8'd234;  #10 
a = 8'd111; b = 8'd235;  #10 
a = 8'd111; b = 8'd236;  #10 
a = 8'd111; b = 8'd237;  #10 
a = 8'd111; b = 8'd238;  #10 
a = 8'd111; b = 8'd239;  #10 
a = 8'd111; b = 8'd240;  #10 
a = 8'd111; b = 8'd241;  #10 
a = 8'd111; b = 8'd242;  #10 
a = 8'd111; b = 8'd243;  #10 
a = 8'd111; b = 8'd244;  #10 
a = 8'd111; b = 8'd245;  #10 
a = 8'd111; b = 8'd246;  #10 
a = 8'd111; b = 8'd247;  #10 
a = 8'd111; b = 8'd248;  #10 
a = 8'd111; b = 8'd249;  #10 
a = 8'd111; b = 8'd250;  #10 
a = 8'd111; b = 8'd251;  #10 
a = 8'd111; b = 8'd252;  #10 
a = 8'd111; b = 8'd253;  #10 
a = 8'd111; b = 8'd254;  #10 
a = 8'd111; b = 8'd255;  #10 
a = 8'd112; b = 8'd0;  #10 
a = 8'd112; b = 8'd1;  #10 
a = 8'd112; b = 8'd2;  #10 
a = 8'd112; b = 8'd3;  #10 
a = 8'd112; b = 8'd4;  #10 
a = 8'd112; b = 8'd5;  #10 
a = 8'd112; b = 8'd6;  #10 
a = 8'd112; b = 8'd7;  #10 
a = 8'd112; b = 8'd8;  #10 
a = 8'd112; b = 8'd9;  #10 
a = 8'd112; b = 8'd10;  #10 
a = 8'd112; b = 8'd11;  #10 
a = 8'd112; b = 8'd12;  #10 
a = 8'd112; b = 8'd13;  #10 
a = 8'd112; b = 8'd14;  #10 
a = 8'd112; b = 8'd15;  #10 
a = 8'd112; b = 8'd16;  #10 
a = 8'd112; b = 8'd17;  #10 
a = 8'd112; b = 8'd18;  #10 
a = 8'd112; b = 8'd19;  #10 
a = 8'd112; b = 8'd20;  #10 
a = 8'd112; b = 8'd21;  #10 
a = 8'd112; b = 8'd22;  #10 
a = 8'd112; b = 8'd23;  #10 
a = 8'd112; b = 8'd24;  #10 
a = 8'd112; b = 8'd25;  #10 
a = 8'd112; b = 8'd26;  #10 
a = 8'd112; b = 8'd27;  #10 
a = 8'd112; b = 8'd28;  #10 
a = 8'd112; b = 8'd29;  #10 
a = 8'd112; b = 8'd30;  #10 
a = 8'd112; b = 8'd31;  #10 
a = 8'd112; b = 8'd32;  #10 
a = 8'd112; b = 8'd33;  #10 
a = 8'd112; b = 8'd34;  #10 
a = 8'd112; b = 8'd35;  #10 
a = 8'd112; b = 8'd36;  #10 
a = 8'd112; b = 8'd37;  #10 
a = 8'd112; b = 8'd38;  #10 
a = 8'd112; b = 8'd39;  #10 
a = 8'd112; b = 8'd40;  #10 
a = 8'd112; b = 8'd41;  #10 
a = 8'd112; b = 8'd42;  #10 
a = 8'd112; b = 8'd43;  #10 
a = 8'd112; b = 8'd44;  #10 
a = 8'd112; b = 8'd45;  #10 
a = 8'd112; b = 8'd46;  #10 
a = 8'd112; b = 8'd47;  #10 
a = 8'd112; b = 8'd48;  #10 
a = 8'd112; b = 8'd49;  #10 
a = 8'd112; b = 8'd50;  #10 
a = 8'd112; b = 8'd51;  #10 
a = 8'd112; b = 8'd52;  #10 
a = 8'd112; b = 8'd53;  #10 
a = 8'd112; b = 8'd54;  #10 
a = 8'd112; b = 8'd55;  #10 
a = 8'd112; b = 8'd56;  #10 
a = 8'd112; b = 8'd57;  #10 
a = 8'd112; b = 8'd58;  #10 
a = 8'd112; b = 8'd59;  #10 
a = 8'd112; b = 8'd60;  #10 
a = 8'd112; b = 8'd61;  #10 
a = 8'd112; b = 8'd62;  #10 
a = 8'd112; b = 8'd63;  #10 
a = 8'd112; b = 8'd64;  #10 
a = 8'd112; b = 8'd65;  #10 
a = 8'd112; b = 8'd66;  #10 
a = 8'd112; b = 8'd67;  #10 
a = 8'd112; b = 8'd68;  #10 
a = 8'd112; b = 8'd69;  #10 
a = 8'd112; b = 8'd70;  #10 
a = 8'd112; b = 8'd71;  #10 
a = 8'd112; b = 8'd72;  #10 
a = 8'd112; b = 8'd73;  #10 
a = 8'd112; b = 8'd74;  #10 
a = 8'd112; b = 8'd75;  #10 
a = 8'd112; b = 8'd76;  #10 
a = 8'd112; b = 8'd77;  #10 
a = 8'd112; b = 8'd78;  #10 
a = 8'd112; b = 8'd79;  #10 
a = 8'd112; b = 8'd80;  #10 
a = 8'd112; b = 8'd81;  #10 
a = 8'd112; b = 8'd82;  #10 
a = 8'd112; b = 8'd83;  #10 
a = 8'd112; b = 8'd84;  #10 
a = 8'd112; b = 8'd85;  #10 
a = 8'd112; b = 8'd86;  #10 
a = 8'd112; b = 8'd87;  #10 
a = 8'd112; b = 8'd88;  #10 
a = 8'd112; b = 8'd89;  #10 
a = 8'd112; b = 8'd90;  #10 
a = 8'd112; b = 8'd91;  #10 
a = 8'd112; b = 8'd92;  #10 
a = 8'd112; b = 8'd93;  #10 
a = 8'd112; b = 8'd94;  #10 
a = 8'd112; b = 8'd95;  #10 
a = 8'd112; b = 8'd96;  #10 
a = 8'd112; b = 8'd97;  #10 
a = 8'd112; b = 8'd98;  #10 
a = 8'd112; b = 8'd99;  #10 
a = 8'd112; b = 8'd100;  #10 
a = 8'd112; b = 8'd101;  #10 
a = 8'd112; b = 8'd102;  #10 
a = 8'd112; b = 8'd103;  #10 
a = 8'd112; b = 8'd104;  #10 
a = 8'd112; b = 8'd105;  #10 
a = 8'd112; b = 8'd106;  #10 
a = 8'd112; b = 8'd107;  #10 
a = 8'd112; b = 8'd108;  #10 
a = 8'd112; b = 8'd109;  #10 
a = 8'd112; b = 8'd110;  #10 
a = 8'd112; b = 8'd111;  #10 
a = 8'd112; b = 8'd112;  #10 
a = 8'd112; b = 8'd113;  #10 
a = 8'd112; b = 8'd114;  #10 
a = 8'd112; b = 8'd115;  #10 
a = 8'd112; b = 8'd116;  #10 
a = 8'd112; b = 8'd117;  #10 
a = 8'd112; b = 8'd118;  #10 
a = 8'd112; b = 8'd119;  #10 
a = 8'd112; b = 8'd120;  #10 
a = 8'd112; b = 8'd121;  #10 
a = 8'd112; b = 8'd122;  #10 
a = 8'd112; b = 8'd123;  #10 
a = 8'd112; b = 8'd124;  #10 
a = 8'd112; b = 8'd125;  #10 
a = 8'd112; b = 8'd126;  #10 
a = 8'd112; b = 8'd127;  #10 
a = 8'd112; b = 8'd128;  #10 
a = 8'd112; b = 8'd129;  #10 
a = 8'd112; b = 8'd130;  #10 
a = 8'd112; b = 8'd131;  #10 
a = 8'd112; b = 8'd132;  #10 
a = 8'd112; b = 8'd133;  #10 
a = 8'd112; b = 8'd134;  #10 
a = 8'd112; b = 8'd135;  #10 
a = 8'd112; b = 8'd136;  #10 
a = 8'd112; b = 8'd137;  #10 
a = 8'd112; b = 8'd138;  #10 
a = 8'd112; b = 8'd139;  #10 
a = 8'd112; b = 8'd140;  #10 
a = 8'd112; b = 8'd141;  #10 
a = 8'd112; b = 8'd142;  #10 
a = 8'd112; b = 8'd143;  #10 
a = 8'd112; b = 8'd144;  #10 
a = 8'd112; b = 8'd145;  #10 
a = 8'd112; b = 8'd146;  #10 
a = 8'd112; b = 8'd147;  #10 
a = 8'd112; b = 8'd148;  #10 
a = 8'd112; b = 8'd149;  #10 
a = 8'd112; b = 8'd150;  #10 
a = 8'd112; b = 8'd151;  #10 
a = 8'd112; b = 8'd152;  #10 
a = 8'd112; b = 8'd153;  #10 
a = 8'd112; b = 8'd154;  #10 
a = 8'd112; b = 8'd155;  #10 
a = 8'd112; b = 8'd156;  #10 
a = 8'd112; b = 8'd157;  #10 
a = 8'd112; b = 8'd158;  #10 
a = 8'd112; b = 8'd159;  #10 
a = 8'd112; b = 8'd160;  #10 
a = 8'd112; b = 8'd161;  #10 
a = 8'd112; b = 8'd162;  #10 
a = 8'd112; b = 8'd163;  #10 
a = 8'd112; b = 8'd164;  #10 
a = 8'd112; b = 8'd165;  #10 
a = 8'd112; b = 8'd166;  #10 
a = 8'd112; b = 8'd167;  #10 
a = 8'd112; b = 8'd168;  #10 
a = 8'd112; b = 8'd169;  #10 
a = 8'd112; b = 8'd170;  #10 
a = 8'd112; b = 8'd171;  #10 
a = 8'd112; b = 8'd172;  #10 
a = 8'd112; b = 8'd173;  #10 
a = 8'd112; b = 8'd174;  #10 
a = 8'd112; b = 8'd175;  #10 
a = 8'd112; b = 8'd176;  #10 
a = 8'd112; b = 8'd177;  #10 
a = 8'd112; b = 8'd178;  #10 
a = 8'd112; b = 8'd179;  #10 
a = 8'd112; b = 8'd180;  #10 
a = 8'd112; b = 8'd181;  #10 
a = 8'd112; b = 8'd182;  #10 
a = 8'd112; b = 8'd183;  #10 
a = 8'd112; b = 8'd184;  #10 
a = 8'd112; b = 8'd185;  #10 
a = 8'd112; b = 8'd186;  #10 
a = 8'd112; b = 8'd187;  #10 
a = 8'd112; b = 8'd188;  #10 
a = 8'd112; b = 8'd189;  #10 
a = 8'd112; b = 8'd190;  #10 
a = 8'd112; b = 8'd191;  #10 
a = 8'd112; b = 8'd192;  #10 
a = 8'd112; b = 8'd193;  #10 
a = 8'd112; b = 8'd194;  #10 
a = 8'd112; b = 8'd195;  #10 
a = 8'd112; b = 8'd196;  #10 
a = 8'd112; b = 8'd197;  #10 
a = 8'd112; b = 8'd198;  #10 
a = 8'd112; b = 8'd199;  #10 
a = 8'd112; b = 8'd200;  #10 
a = 8'd112; b = 8'd201;  #10 
a = 8'd112; b = 8'd202;  #10 
a = 8'd112; b = 8'd203;  #10 
a = 8'd112; b = 8'd204;  #10 
a = 8'd112; b = 8'd205;  #10 
a = 8'd112; b = 8'd206;  #10 
a = 8'd112; b = 8'd207;  #10 
a = 8'd112; b = 8'd208;  #10 
a = 8'd112; b = 8'd209;  #10 
a = 8'd112; b = 8'd210;  #10 
a = 8'd112; b = 8'd211;  #10 
a = 8'd112; b = 8'd212;  #10 
a = 8'd112; b = 8'd213;  #10 
a = 8'd112; b = 8'd214;  #10 
a = 8'd112; b = 8'd215;  #10 
a = 8'd112; b = 8'd216;  #10 
a = 8'd112; b = 8'd217;  #10 
a = 8'd112; b = 8'd218;  #10 
a = 8'd112; b = 8'd219;  #10 
a = 8'd112; b = 8'd220;  #10 
a = 8'd112; b = 8'd221;  #10 
a = 8'd112; b = 8'd222;  #10 
a = 8'd112; b = 8'd223;  #10 
a = 8'd112; b = 8'd224;  #10 
a = 8'd112; b = 8'd225;  #10 
a = 8'd112; b = 8'd226;  #10 
a = 8'd112; b = 8'd227;  #10 
a = 8'd112; b = 8'd228;  #10 
a = 8'd112; b = 8'd229;  #10 
a = 8'd112; b = 8'd230;  #10 
a = 8'd112; b = 8'd231;  #10 
a = 8'd112; b = 8'd232;  #10 
a = 8'd112; b = 8'd233;  #10 
a = 8'd112; b = 8'd234;  #10 
a = 8'd112; b = 8'd235;  #10 
a = 8'd112; b = 8'd236;  #10 
a = 8'd112; b = 8'd237;  #10 
a = 8'd112; b = 8'd238;  #10 
a = 8'd112; b = 8'd239;  #10 
a = 8'd112; b = 8'd240;  #10 
a = 8'd112; b = 8'd241;  #10 
a = 8'd112; b = 8'd242;  #10 
a = 8'd112; b = 8'd243;  #10 
a = 8'd112; b = 8'd244;  #10 
a = 8'd112; b = 8'd245;  #10 
a = 8'd112; b = 8'd246;  #10 
a = 8'd112; b = 8'd247;  #10 
a = 8'd112; b = 8'd248;  #10 
a = 8'd112; b = 8'd249;  #10 
a = 8'd112; b = 8'd250;  #10 
a = 8'd112; b = 8'd251;  #10 
a = 8'd112; b = 8'd252;  #10 
a = 8'd112; b = 8'd253;  #10 
a = 8'd112; b = 8'd254;  #10 
a = 8'd112; b = 8'd255;  #10 
a = 8'd113; b = 8'd0;  #10 
a = 8'd113; b = 8'd1;  #10 
a = 8'd113; b = 8'd2;  #10 
a = 8'd113; b = 8'd3;  #10 
a = 8'd113; b = 8'd4;  #10 
a = 8'd113; b = 8'd5;  #10 
a = 8'd113; b = 8'd6;  #10 
a = 8'd113; b = 8'd7;  #10 
a = 8'd113; b = 8'd8;  #10 
a = 8'd113; b = 8'd9;  #10 
a = 8'd113; b = 8'd10;  #10 
a = 8'd113; b = 8'd11;  #10 
a = 8'd113; b = 8'd12;  #10 
a = 8'd113; b = 8'd13;  #10 
a = 8'd113; b = 8'd14;  #10 
a = 8'd113; b = 8'd15;  #10 
a = 8'd113; b = 8'd16;  #10 
a = 8'd113; b = 8'd17;  #10 
a = 8'd113; b = 8'd18;  #10 
a = 8'd113; b = 8'd19;  #10 
a = 8'd113; b = 8'd20;  #10 
a = 8'd113; b = 8'd21;  #10 
a = 8'd113; b = 8'd22;  #10 
a = 8'd113; b = 8'd23;  #10 
a = 8'd113; b = 8'd24;  #10 
a = 8'd113; b = 8'd25;  #10 
a = 8'd113; b = 8'd26;  #10 
a = 8'd113; b = 8'd27;  #10 
a = 8'd113; b = 8'd28;  #10 
a = 8'd113; b = 8'd29;  #10 
a = 8'd113; b = 8'd30;  #10 
a = 8'd113; b = 8'd31;  #10 
a = 8'd113; b = 8'd32;  #10 
a = 8'd113; b = 8'd33;  #10 
a = 8'd113; b = 8'd34;  #10 
a = 8'd113; b = 8'd35;  #10 
a = 8'd113; b = 8'd36;  #10 
a = 8'd113; b = 8'd37;  #10 
a = 8'd113; b = 8'd38;  #10 
a = 8'd113; b = 8'd39;  #10 
a = 8'd113; b = 8'd40;  #10 
a = 8'd113; b = 8'd41;  #10 
a = 8'd113; b = 8'd42;  #10 
a = 8'd113; b = 8'd43;  #10 
a = 8'd113; b = 8'd44;  #10 
a = 8'd113; b = 8'd45;  #10 
a = 8'd113; b = 8'd46;  #10 
a = 8'd113; b = 8'd47;  #10 
a = 8'd113; b = 8'd48;  #10 
a = 8'd113; b = 8'd49;  #10 
a = 8'd113; b = 8'd50;  #10 
a = 8'd113; b = 8'd51;  #10 
a = 8'd113; b = 8'd52;  #10 
a = 8'd113; b = 8'd53;  #10 
a = 8'd113; b = 8'd54;  #10 
a = 8'd113; b = 8'd55;  #10 
a = 8'd113; b = 8'd56;  #10 
a = 8'd113; b = 8'd57;  #10 
a = 8'd113; b = 8'd58;  #10 
a = 8'd113; b = 8'd59;  #10 
a = 8'd113; b = 8'd60;  #10 
a = 8'd113; b = 8'd61;  #10 
a = 8'd113; b = 8'd62;  #10 
a = 8'd113; b = 8'd63;  #10 
a = 8'd113; b = 8'd64;  #10 
a = 8'd113; b = 8'd65;  #10 
a = 8'd113; b = 8'd66;  #10 
a = 8'd113; b = 8'd67;  #10 
a = 8'd113; b = 8'd68;  #10 
a = 8'd113; b = 8'd69;  #10 
a = 8'd113; b = 8'd70;  #10 
a = 8'd113; b = 8'd71;  #10 
a = 8'd113; b = 8'd72;  #10 
a = 8'd113; b = 8'd73;  #10 
a = 8'd113; b = 8'd74;  #10 
a = 8'd113; b = 8'd75;  #10 
a = 8'd113; b = 8'd76;  #10 
a = 8'd113; b = 8'd77;  #10 
a = 8'd113; b = 8'd78;  #10 
a = 8'd113; b = 8'd79;  #10 
a = 8'd113; b = 8'd80;  #10 
a = 8'd113; b = 8'd81;  #10 
a = 8'd113; b = 8'd82;  #10 
a = 8'd113; b = 8'd83;  #10 
a = 8'd113; b = 8'd84;  #10 
a = 8'd113; b = 8'd85;  #10 
a = 8'd113; b = 8'd86;  #10 
a = 8'd113; b = 8'd87;  #10 
a = 8'd113; b = 8'd88;  #10 
a = 8'd113; b = 8'd89;  #10 
a = 8'd113; b = 8'd90;  #10 
a = 8'd113; b = 8'd91;  #10 
a = 8'd113; b = 8'd92;  #10 
a = 8'd113; b = 8'd93;  #10 
a = 8'd113; b = 8'd94;  #10 
a = 8'd113; b = 8'd95;  #10 
a = 8'd113; b = 8'd96;  #10 
a = 8'd113; b = 8'd97;  #10 
a = 8'd113; b = 8'd98;  #10 
a = 8'd113; b = 8'd99;  #10 
a = 8'd113; b = 8'd100;  #10 
a = 8'd113; b = 8'd101;  #10 
a = 8'd113; b = 8'd102;  #10 
a = 8'd113; b = 8'd103;  #10 
a = 8'd113; b = 8'd104;  #10 
a = 8'd113; b = 8'd105;  #10 
a = 8'd113; b = 8'd106;  #10 
a = 8'd113; b = 8'd107;  #10 
a = 8'd113; b = 8'd108;  #10 
a = 8'd113; b = 8'd109;  #10 
a = 8'd113; b = 8'd110;  #10 
a = 8'd113; b = 8'd111;  #10 
a = 8'd113; b = 8'd112;  #10 
a = 8'd113; b = 8'd113;  #10 
a = 8'd113; b = 8'd114;  #10 
a = 8'd113; b = 8'd115;  #10 
a = 8'd113; b = 8'd116;  #10 
a = 8'd113; b = 8'd117;  #10 
a = 8'd113; b = 8'd118;  #10 
a = 8'd113; b = 8'd119;  #10 
a = 8'd113; b = 8'd120;  #10 
a = 8'd113; b = 8'd121;  #10 
a = 8'd113; b = 8'd122;  #10 
a = 8'd113; b = 8'd123;  #10 
a = 8'd113; b = 8'd124;  #10 
a = 8'd113; b = 8'd125;  #10 
a = 8'd113; b = 8'd126;  #10 
a = 8'd113; b = 8'd127;  #10 
a = 8'd113; b = 8'd128;  #10 
a = 8'd113; b = 8'd129;  #10 
a = 8'd113; b = 8'd130;  #10 
a = 8'd113; b = 8'd131;  #10 
a = 8'd113; b = 8'd132;  #10 
a = 8'd113; b = 8'd133;  #10 
a = 8'd113; b = 8'd134;  #10 
a = 8'd113; b = 8'd135;  #10 
a = 8'd113; b = 8'd136;  #10 
a = 8'd113; b = 8'd137;  #10 
a = 8'd113; b = 8'd138;  #10 
a = 8'd113; b = 8'd139;  #10 
a = 8'd113; b = 8'd140;  #10 
a = 8'd113; b = 8'd141;  #10 
a = 8'd113; b = 8'd142;  #10 
a = 8'd113; b = 8'd143;  #10 
a = 8'd113; b = 8'd144;  #10 
a = 8'd113; b = 8'd145;  #10 
a = 8'd113; b = 8'd146;  #10 
a = 8'd113; b = 8'd147;  #10 
a = 8'd113; b = 8'd148;  #10 
a = 8'd113; b = 8'd149;  #10 
a = 8'd113; b = 8'd150;  #10 
a = 8'd113; b = 8'd151;  #10 
a = 8'd113; b = 8'd152;  #10 
a = 8'd113; b = 8'd153;  #10 
a = 8'd113; b = 8'd154;  #10 
a = 8'd113; b = 8'd155;  #10 
a = 8'd113; b = 8'd156;  #10 
a = 8'd113; b = 8'd157;  #10 
a = 8'd113; b = 8'd158;  #10 
a = 8'd113; b = 8'd159;  #10 
a = 8'd113; b = 8'd160;  #10 
a = 8'd113; b = 8'd161;  #10 
a = 8'd113; b = 8'd162;  #10 
a = 8'd113; b = 8'd163;  #10 
a = 8'd113; b = 8'd164;  #10 
a = 8'd113; b = 8'd165;  #10 
a = 8'd113; b = 8'd166;  #10 
a = 8'd113; b = 8'd167;  #10 
a = 8'd113; b = 8'd168;  #10 
a = 8'd113; b = 8'd169;  #10 
a = 8'd113; b = 8'd170;  #10 
a = 8'd113; b = 8'd171;  #10 
a = 8'd113; b = 8'd172;  #10 
a = 8'd113; b = 8'd173;  #10 
a = 8'd113; b = 8'd174;  #10 
a = 8'd113; b = 8'd175;  #10 
a = 8'd113; b = 8'd176;  #10 
a = 8'd113; b = 8'd177;  #10 
a = 8'd113; b = 8'd178;  #10 
a = 8'd113; b = 8'd179;  #10 
a = 8'd113; b = 8'd180;  #10 
a = 8'd113; b = 8'd181;  #10 
a = 8'd113; b = 8'd182;  #10 
a = 8'd113; b = 8'd183;  #10 
a = 8'd113; b = 8'd184;  #10 
a = 8'd113; b = 8'd185;  #10 
a = 8'd113; b = 8'd186;  #10 
a = 8'd113; b = 8'd187;  #10 
a = 8'd113; b = 8'd188;  #10 
a = 8'd113; b = 8'd189;  #10 
a = 8'd113; b = 8'd190;  #10 
a = 8'd113; b = 8'd191;  #10 
a = 8'd113; b = 8'd192;  #10 
a = 8'd113; b = 8'd193;  #10 
a = 8'd113; b = 8'd194;  #10 
a = 8'd113; b = 8'd195;  #10 
a = 8'd113; b = 8'd196;  #10 
a = 8'd113; b = 8'd197;  #10 
a = 8'd113; b = 8'd198;  #10 
a = 8'd113; b = 8'd199;  #10 
a = 8'd113; b = 8'd200;  #10 
a = 8'd113; b = 8'd201;  #10 
a = 8'd113; b = 8'd202;  #10 
a = 8'd113; b = 8'd203;  #10 
a = 8'd113; b = 8'd204;  #10 
a = 8'd113; b = 8'd205;  #10 
a = 8'd113; b = 8'd206;  #10 
a = 8'd113; b = 8'd207;  #10 
a = 8'd113; b = 8'd208;  #10 
a = 8'd113; b = 8'd209;  #10 
a = 8'd113; b = 8'd210;  #10 
a = 8'd113; b = 8'd211;  #10 
a = 8'd113; b = 8'd212;  #10 
a = 8'd113; b = 8'd213;  #10 
a = 8'd113; b = 8'd214;  #10 
a = 8'd113; b = 8'd215;  #10 
a = 8'd113; b = 8'd216;  #10 
a = 8'd113; b = 8'd217;  #10 
a = 8'd113; b = 8'd218;  #10 
a = 8'd113; b = 8'd219;  #10 
a = 8'd113; b = 8'd220;  #10 
a = 8'd113; b = 8'd221;  #10 
a = 8'd113; b = 8'd222;  #10 
a = 8'd113; b = 8'd223;  #10 
a = 8'd113; b = 8'd224;  #10 
a = 8'd113; b = 8'd225;  #10 
a = 8'd113; b = 8'd226;  #10 
a = 8'd113; b = 8'd227;  #10 
a = 8'd113; b = 8'd228;  #10 
a = 8'd113; b = 8'd229;  #10 
a = 8'd113; b = 8'd230;  #10 
a = 8'd113; b = 8'd231;  #10 
a = 8'd113; b = 8'd232;  #10 
a = 8'd113; b = 8'd233;  #10 
a = 8'd113; b = 8'd234;  #10 
a = 8'd113; b = 8'd235;  #10 
a = 8'd113; b = 8'd236;  #10 
a = 8'd113; b = 8'd237;  #10 
a = 8'd113; b = 8'd238;  #10 
a = 8'd113; b = 8'd239;  #10 
a = 8'd113; b = 8'd240;  #10 
a = 8'd113; b = 8'd241;  #10 
a = 8'd113; b = 8'd242;  #10 
a = 8'd113; b = 8'd243;  #10 
a = 8'd113; b = 8'd244;  #10 
a = 8'd113; b = 8'd245;  #10 
a = 8'd113; b = 8'd246;  #10 
a = 8'd113; b = 8'd247;  #10 
a = 8'd113; b = 8'd248;  #10 
a = 8'd113; b = 8'd249;  #10 
a = 8'd113; b = 8'd250;  #10 
a = 8'd113; b = 8'd251;  #10 
a = 8'd113; b = 8'd252;  #10 
a = 8'd113; b = 8'd253;  #10 
a = 8'd113; b = 8'd254;  #10 
a = 8'd113; b = 8'd255;  #10 
a = 8'd114; b = 8'd0;  #10 
a = 8'd114; b = 8'd1;  #10 
a = 8'd114; b = 8'd2;  #10 
a = 8'd114; b = 8'd3;  #10 
a = 8'd114; b = 8'd4;  #10 
a = 8'd114; b = 8'd5;  #10 
a = 8'd114; b = 8'd6;  #10 
a = 8'd114; b = 8'd7;  #10 
a = 8'd114; b = 8'd8;  #10 
a = 8'd114; b = 8'd9;  #10 
a = 8'd114; b = 8'd10;  #10 
a = 8'd114; b = 8'd11;  #10 
a = 8'd114; b = 8'd12;  #10 
a = 8'd114; b = 8'd13;  #10 
a = 8'd114; b = 8'd14;  #10 
a = 8'd114; b = 8'd15;  #10 
a = 8'd114; b = 8'd16;  #10 
a = 8'd114; b = 8'd17;  #10 
a = 8'd114; b = 8'd18;  #10 
a = 8'd114; b = 8'd19;  #10 
a = 8'd114; b = 8'd20;  #10 
a = 8'd114; b = 8'd21;  #10 
a = 8'd114; b = 8'd22;  #10 
a = 8'd114; b = 8'd23;  #10 
a = 8'd114; b = 8'd24;  #10 
a = 8'd114; b = 8'd25;  #10 
a = 8'd114; b = 8'd26;  #10 
a = 8'd114; b = 8'd27;  #10 
a = 8'd114; b = 8'd28;  #10 
a = 8'd114; b = 8'd29;  #10 
a = 8'd114; b = 8'd30;  #10 
a = 8'd114; b = 8'd31;  #10 
a = 8'd114; b = 8'd32;  #10 
a = 8'd114; b = 8'd33;  #10 
a = 8'd114; b = 8'd34;  #10 
a = 8'd114; b = 8'd35;  #10 
a = 8'd114; b = 8'd36;  #10 
a = 8'd114; b = 8'd37;  #10 
a = 8'd114; b = 8'd38;  #10 
a = 8'd114; b = 8'd39;  #10 
a = 8'd114; b = 8'd40;  #10 
a = 8'd114; b = 8'd41;  #10 
a = 8'd114; b = 8'd42;  #10 
a = 8'd114; b = 8'd43;  #10 
a = 8'd114; b = 8'd44;  #10 
a = 8'd114; b = 8'd45;  #10 
a = 8'd114; b = 8'd46;  #10 
a = 8'd114; b = 8'd47;  #10 
a = 8'd114; b = 8'd48;  #10 
a = 8'd114; b = 8'd49;  #10 
a = 8'd114; b = 8'd50;  #10 
a = 8'd114; b = 8'd51;  #10 
a = 8'd114; b = 8'd52;  #10 
a = 8'd114; b = 8'd53;  #10 
a = 8'd114; b = 8'd54;  #10 
a = 8'd114; b = 8'd55;  #10 
a = 8'd114; b = 8'd56;  #10 
a = 8'd114; b = 8'd57;  #10 
a = 8'd114; b = 8'd58;  #10 
a = 8'd114; b = 8'd59;  #10 
a = 8'd114; b = 8'd60;  #10 
a = 8'd114; b = 8'd61;  #10 
a = 8'd114; b = 8'd62;  #10 
a = 8'd114; b = 8'd63;  #10 
a = 8'd114; b = 8'd64;  #10 
a = 8'd114; b = 8'd65;  #10 
a = 8'd114; b = 8'd66;  #10 
a = 8'd114; b = 8'd67;  #10 
a = 8'd114; b = 8'd68;  #10 
a = 8'd114; b = 8'd69;  #10 
a = 8'd114; b = 8'd70;  #10 
a = 8'd114; b = 8'd71;  #10 
a = 8'd114; b = 8'd72;  #10 
a = 8'd114; b = 8'd73;  #10 
a = 8'd114; b = 8'd74;  #10 
a = 8'd114; b = 8'd75;  #10 
a = 8'd114; b = 8'd76;  #10 
a = 8'd114; b = 8'd77;  #10 
a = 8'd114; b = 8'd78;  #10 
a = 8'd114; b = 8'd79;  #10 
a = 8'd114; b = 8'd80;  #10 
a = 8'd114; b = 8'd81;  #10 
a = 8'd114; b = 8'd82;  #10 
a = 8'd114; b = 8'd83;  #10 
a = 8'd114; b = 8'd84;  #10 
a = 8'd114; b = 8'd85;  #10 
a = 8'd114; b = 8'd86;  #10 
a = 8'd114; b = 8'd87;  #10 
a = 8'd114; b = 8'd88;  #10 
a = 8'd114; b = 8'd89;  #10 
a = 8'd114; b = 8'd90;  #10 
a = 8'd114; b = 8'd91;  #10 
a = 8'd114; b = 8'd92;  #10 
a = 8'd114; b = 8'd93;  #10 
a = 8'd114; b = 8'd94;  #10 
a = 8'd114; b = 8'd95;  #10 
a = 8'd114; b = 8'd96;  #10 
a = 8'd114; b = 8'd97;  #10 
a = 8'd114; b = 8'd98;  #10 
a = 8'd114; b = 8'd99;  #10 
a = 8'd114; b = 8'd100;  #10 
a = 8'd114; b = 8'd101;  #10 
a = 8'd114; b = 8'd102;  #10 
a = 8'd114; b = 8'd103;  #10 
a = 8'd114; b = 8'd104;  #10 
a = 8'd114; b = 8'd105;  #10 
a = 8'd114; b = 8'd106;  #10 
a = 8'd114; b = 8'd107;  #10 
a = 8'd114; b = 8'd108;  #10 
a = 8'd114; b = 8'd109;  #10 
a = 8'd114; b = 8'd110;  #10 
a = 8'd114; b = 8'd111;  #10 
a = 8'd114; b = 8'd112;  #10 
a = 8'd114; b = 8'd113;  #10 
a = 8'd114; b = 8'd114;  #10 
a = 8'd114; b = 8'd115;  #10 
a = 8'd114; b = 8'd116;  #10 
a = 8'd114; b = 8'd117;  #10 
a = 8'd114; b = 8'd118;  #10 
a = 8'd114; b = 8'd119;  #10 
a = 8'd114; b = 8'd120;  #10 
a = 8'd114; b = 8'd121;  #10 
a = 8'd114; b = 8'd122;  #10 
a = 8'd114; b = 8'd123;  #10 
a = 8'd114; b = 8'd124;  #10 
a = 8'd114; b = 8'd125;  #10 
a = 8'd114; b = 8'd126;  #10 
a = 8'd114; b = 8'd127;  #10 
a = 8'd114; b = 8'd128;  #10 
a = 8'd114; b = 8'd129;  #10 
a = 8'd114; b = 8'd130;  #10 
a = 8'd114; b = 8'd131;  #10 
a = 8'd114; b = 8'd132;  #10 
a = 8'd114; b = 8'd133;  #10 
a = 8'd114; b = 8'd134;  #10 
a = 8'd114; b = 8'd135;  #10 
a = 8'd114; b = 8'd136;  #10 
a = 8'd114; b = 8'd137;  #10 
a = 8'd114; b = 8'd138;  #10 
a = 8'd114; b = 8'd139;  #10 
a = 8'd114; b = 8'd140;  #10 
a = 8'd114; b = 8'd141;  #10 
a = 8'd114; b = 8'd142;  #10 
a = 8'd114; b = 8'd143;  #10 
a = 8'd114; b = 8'd144;  #10 
a = 8'd114; b = 8'd145;  #10 
a = 8'd114; b = 8'd146;  #10 
a = 8'd114; b = 8'd147;  #10 
a = 8'd114; b = 8'd148;  #10 
a = 8'd114; b = 8'd149;  #10 
a = 8'd114; b = 8'd150;  #10 
a = 8'd114; b = 8'd151;  #10 
a = 8'd114; b = 8'd152;  #10 
a = 8'd114; b = 8'd153;  #10 
a = 8'd114; b = 8'd154;  #10 
a = 8'd114; b = 8'd155;  #10 
a = 8'd114; b = 8'd156;  #10 
a = 8'd114; b = 8'd157;  #10 
a = 8'd114; b = 8'd158;  #10 
a = 8'd114; b = 8'd159;  #10 
a = 8'd114; b = 8'd160;  #10 
a = 8'd114; b = 8'd161;  #10 
a = 8'd114; b = 8'd162;  #10 
a = 8'd114; b = 8'd163;  #10 
a = 8'd114; b = 8'd164;  #10 
a = 8'd114; b = 8'd165;  #10 
a = 8'd114; b = 8'd166;  #10 
a = 8'd114; b = 8'd167;  #10 
a = 8'd114; b = 8'd168;  #10 
a = 8'd114; b = 8'd169;  #10 
a = 8'd114; b = 8'd170;  #10 
a = 8'd114; b = 8'd171;  #10 
a = 8'd114; b = 8'd172;  #10 
a = 8'd114; b = 8'd173;  #10 
a = 8'd114; b = 8'd174;  #10 
a = 8'd114; b = 8'd175;  #10 
a = 8'd114; b = 8'd176;  #10 
a = 8'd114; b = 8'd177;  #10 
a = 8'd114; b = 8'd178;  #10 
a = 8'd114; b = 8'd179;  #10 
a = 8'd114; b = 8'd180;  #10 
a = 8'd114; b = 8'd181;  #10 
a = 8'd114; b = 8'd182;  #10 
a = 8'd114; b = 8'd183;  #10 
a = 8'd114; b = 8'd184;  #10 
a = 8'd114; b = 8'd185;  #10 
a = 8'd114; b = 8'd186;  #10 
a = 8'd114; b = 8'd187;  #10 
a = 8'd114; b = 8'd188;  #10 
a = 8'd114; b = 8'd189;  #10 
a = 8'd114; b = 8'd190;  #10 
a = 8'd114; b = 8'd191;  #10 
a = 8'd114; b = 8'd192;  #10 
a = 8'd114; b = 8'd193;  #10 
a = 8'd114; b = 8'd194;  #10 
a = 8'd114; b = 8'd195;  #10 
a = 8'd114; b = 8'd196;  #10 
a = 8'd114; b = 8'd197;  #10 
a = 8'd114; b = 8'd198;  #10 
a = 8'd114; b = 8'd199;  #10 
a = 8'd114; b = 8'd200;  #10 
a = 8'd114; b = 8'd201;  #10 
a = 8'd114; b = 8'd202;  #10 
a = 8'd114; b = 8'd203;  #10 
a = 8'd114; b = 8'd204;  #10 
a = 8'd114; b = 8'd205;  #10 
a = 8'd114; b = 8'd206;  #10 
a = 8'd114; b = 8'd207;  #10 
a = 8'd114; b = 8'd208;  #10 
a = 8'd114; b = 8'd209;  #10 
a = 8'd114; b = 8'd210;  #10 
a = 8'd114; b = 8'd211;  #10 
a = 8'd114; b = 8'd212;  #10 
a = 8'd114; b = 8'd213;  #10 
a = 8'd114; b = 8'd214;  #10 
a = 8'd114; b = 8'd215;  #10 
a = 8'd114; b = 8'd216;  #10 
a = 8'd114; b = 8'd217;  #10 
a = 8'd114; b = 8'd218;  #10 
a = 8'd114; b = 8'd219;  #10 
a = 8'd114; b = 8'd220;  #10 
a = 8'd114; b = 8'd221;  #10 
a = 8'd114; b = 8'd222;  #10 
a = 8'd114; b = 8'd223;  #10 
a = 8'd114; b = 8'd224;  #10 
a = 8'd114; b = 8'd225;  #10 
a = 8'd114; b = 8'd226;  #10 
a = 8'd114; b = 8'd227;  #10 
a = 8'd114; b = 8'd228;  #10 
a = 8'd114; b = 8'd229;  #10 
a = 8'd114; b = 8'd230;  #10 
a = 8'd114; b = 8'd231;  #10 
a = 8'd114; b = 8'd232;  #10 
a = 8'd114; b = 8'd233;  #10 
a = 8'd114; b = 8'd234;  #10 
a = 8'd114; b = 8'd235;  #10 
a = 8'd114; b = 8'd236;  #10 
a = 8'd114; b = 8'd237;  #10 
a = 8'd114; b = 8'd238;  #10 
a = 8'd114; b = 8'd239;  #10 
a = 8'd114; b = 8'd240;  #10 
a = 8'd114; b = 8'd241;  #10 
a = 8'd114; b = 8'd242;  #10 
a = 8'd114; b = 8'd243;  #10 
a = 8'd114; b = 8'd244;  #10 
a = 8'd114; b = 8'd245;  #10 
a = 8'd114; b = 8'd246;  #10 
a = 8'd114; b = 8'd247;  #10 
a = 8'd114; b = 8'd248;  #10 
a = 8'd114; b = 8'd249;  #10 
a = 8'd114; b = 8'd250;  #10 
a = 8'd114; b = 8'd251;  #10 
a = 8'd114; b = 8'd252;  #10 
a = 8'd114; b = 8'd253;  #10 
a = 8'd114; b = 8'd254;  #10 
a = 8'd114; b = 8'd255;  #10 
a = 8'd115; b = 8'd0;  #10 
a = 8'd115; b = 8'd1;  #10 
a = 8'd115; b = 8'd2;  #10 
a = 8'd115; b = 8'd3;  #10 
a = 8'd115; b = 8'd4;  #10 
a = 8'd115; b = 8'd5;  #10 
a = 8'd115; b = 8'd6;  #10 
a = 8'd115; b = 8'd7;  #10 
a = 8'd115; b = 8'd8;  #10 
a = 8'd115; b = 8'd9;  #10 
a = 8'd115; b = 8'd10;  #10 
a = 8'd115; b = 8'd11;  #10 
a = 8'd115; b = 8'd12;  #10 
a = 8'd115; b = 8'd13;  #10 
a = 8'd115; b = 8'd14;  #10 
a = 8'd115; b = 8'd15;  #10 
a = 8'd115; b = 8'd16;  #10 
a = 8'd115; b = 8'd17;  #10 
a = 8'd115; b = 8'd18;  #10 
a = 8'd115; b = 8'd19;  #10 
a = 8'd115; b = 8'd20;  #10 
a = 8'd115; b = 8'd21;  #10 
a = 8'd115; b = 8'd22;  #10 
a = 8'd115; b = 8'd23;  #10 
a = 8'd115; b = 8'd24;  #10 
a = 8'd115; b = 8'd25;  #10 
a = 8'd115; b = 8'd26;  #10 
a = 8'd115; b = 8'd27;  #10 
a = 8'd115; b = 8'd28;  #10 
a = 8'd115; b = 8'd29;  #10 
a = 8'd115; b = 8'd30;  #10 
a = 8'd115; b = 8'd31;  #10 
a = 8'd115; b = 8'd32;  #10 
a = 8'd115; b = 8'd33;  #10 
a = 8'd115; b = 8'd34;  #10 
a = 8'd115; b = 8'd35;  #10 
a = 8'd115; b = 8'd36;  #10 
a = 8'd115; b = 8'd37;  #10 
a = 8'd115; b = 8'd38;  #10 
a = 8'd115; b = 8'd39;  #10 
a = 8'd115; b = 8'd40;  #10 
a = 8'd115; b = 8'd41;  #10 
a = 8'd115; b = 8'd42;  #10 
a = 8'd115; b = 8'd43;  #10 
a = 8'd115; b = 8'd44;  #10 
a = 8'd115; b = 8'd45;  #10 
a = 8'd115; b = 8'd46;  #10 
a = 8'd115; b = 8'd47;  #10 
a = 8'd115; b = 8'd48;  #10 
a = 8'd115; b = 8'd49;  #10 
a = 8'd115; b = 8'd50;  #10 
a = 8'd115; b = 8'd51;  #10 
a = 8'd115; b = 8'd52;  #10 
a = 8'd115; b = 8'd53;  #10 
a = 8'd115; b = 8'd54;  #10 
a = 8'd115; b = 8'd55;  #10 
a = 8'd115; b = 8'd56;  #10 
a = 8'd115; b = 8'd57;  #10 
a = 8'd115; b = 8'd58;  #10 
a = 8'd115; b = 8'd59;  #10 
a = 8'd115; b = 8'd60;  #10 
a = 8'd115; b = 8'd61;  #10 
a = 8'd115; b = 8'd62;  #10 
a = 8'd115; b = 8'd63;  #10 
a = 8'd115; b = 8'd64;  #10 
a = 8'd115; b = 8'd65;  #10 
a = 8'd115; b = 8'd66;  #10 
a = 8'd115; b = 8'd67;  #10 
a = 8'd115; b = 8'd68;  #10 
a = 8'd115; b = 8'd69;  #10 
a = 8'd115; b = 8'd70;  #10 
a = 8'd115; b = 8'd71;  #10 
a = 8'd115; b = 8'd72;  #10 
a = 8'd115; b = 8'd73;  #10 
a = 8'd115; b = 8'd74;  #10 
a = 8'd115; b = 8'd75;  #10 
a = 8'd115; b = 8'd76;  #10 
a = 8'd115; b = 8'd77;  #10 
a = 8'd115; b = 8'd78;  #10 
a = 8'd115; b = 8'd79;  #10 
a = 8'd115; b = 8'd80;  #10 
a = 8'd115; b = 8'd81;  #10 
a = 8'd115; b = 8'd82;  #10 
a = 8'd115; b = 8'd83;  #10 
a = 8'd115; b = 8'd84;  #10 
a = 8'd115; b = 8'd85;  #10 
a = 8'd115; b = 8'd86;  #10 
a = 8'd115; b = 8'd87;  #10 
a = 8'd115; b = 8'd88;  #10 
a = 8'd115; b = 8'd89;  #10 
a = 8'd115; b = 8'd90;  #10 
a = 8'd115; b = 8'd91;  #10 
a = 8'd115; b = 8'd92;  #10 
a = 8'd115; b = 8'd93;  #10 
a = 8'd115; b = 8'd94;  #10 
a = 8'd115; b = 8'd95;  #10 
a = 8'd115; b = 8'd96;  #10 
a = 8'd115; b = 8'd97;  #10 
a = 8'd115; b = 8'd98;  #10 
a = 8'd115; b = 8'd99;  #10 
a = 8'd115; b = 8'd100;  #10 
a = 8'd115; b = 8'd101;  #10 
a = 8'd115; b = 8'd102;  #10 
a = 8'd115; b = 8'd103;  #10 
a = 8'd115; b = 8'd104;  #10 
a = 8'd115; b = 8'd105;  #10 
a = 8'd115; b = 8'd106;  #10 
a = 8'd115; b = 8'd107;  #10 
a = 8'd115; b = 8'd108;  #10 
a = 8'd115; b = 8'd109;  #10 
a = 8'd115; b = 8'd110;  #10 
a = 8'd115; b = 8'd111;  #10 
a = 8'd115; b = 8'd112;  #10 
a = 8'd115; b = 8'd113;  #10 
a = 8'd115; b = 8'd114;  #10 
a = 8'd115; b = 8'd115;  #10 
a = 8'd115; b = 8'd116;  #10 
a = 8'd115; b = 8'd117;  #10 
a = 8'd115; b = 8'd118;  #10 
a = 8'd115; b = 8'd119;  #10 
a = 8'd115; b = 8'd120;  #10 
a = 8'd115; b = 8'd121;  #10 
a = 8'd115; b = 8'd122;  #10 
a = 8'd115; b = 8'd123;  #10 
a = 8'd115; b = 8'd124;  #10 
a = 8'd115; b = 8'd125;  #10 
a = 8'd115; b = 8'd126;  #10 
a = 8'd115; b = 8'd127;  #10 
a = 8'd115; b = 8'd128;  #10 
a = 8'd115; b = 8'd129;  #10 
a = 8'd115; b = 8'd130;  #10 
a = 8'd115; b = 8'd131;  #10 
a = 8'd115; b = 8'd132;  #10 
a = 8'd115; b = 8'd133;  #10 
a = 8'd115; b = 8'd134;  #10 
a = 8'd115; b = 8'd135;  #10 
a = 8'd115; b = 8'd136;  #10 
a = 8'd115; b = 8'd137;  #10 
a = 8'd115; b = 8'd138;  #10 
a = 8'd115; b = 8'd139;  #10 
a = 8'd115; b = 8'd140;  #10 
a = 8'd115; b = 8'd141;  #10 
a = 8'd115; b = 8'd142;  #10 
a = 8'd115; b = 8'd143;  #10 
a = 8'd115; b = 8'd144;  #10 
a = 8'd115; b = 8'd145;  #10 
a = 8'd115; b = 8'd146;  #10 
a = 8'd115; b = 8'd147;  #10 
a = 8'd115; b = 8'd148;  #10 
a = 8'd115; b = 8'd149;  #10 
a = 8'd115; b = 8'd150;  #10 
a = 8'd115; b = 8'd151;  #10 
a = 8'd115; b = 8'd152;  #10 
a = 8'd115; b = 8'd153;  #10 
a = 8'd115; b = 8'd154;  #10 
a = 8'd115; b = 8'd155;  #10 
a = 8'd115; b = 8'd156;  #10 
a = 8'd115; b = 8'd157;  #10 
a = 8'd115; b = 8'd158;  #10 
a = 8'd115; b = 8'd159;  #10 
a = 8'd115; b = 8'd160;  #10 
a = 8'd115; b = 8'd161;  #10 
a = 8'd115; b = 8'd162;  #10 
a = 8'd115; b = 8'd163;  #10 
a = 8'd115; b = 8'd164;  #10 
a = 8'd115; b = 8'd165;  #10 
a = 8'd115; b = 8'd166;  #10 
a = 8'd115; b = 8'd167;  #10 
a = 8'd115; b = 8'd168;  #10 
a = 8'd115; b = 8'd169;  #10 
a = 8'd115; b = 8'd170;  #10 
a = 8'd115; b = 8'd171;  #10 
a = 8'd115; b = 8'd172;  #10 
a = 8'd115; b = 8'd173;  #10 
a = 8'd115; b = 8'd174;  #10 
a = 8'd115; b = 8'd175;  #10 
a = 8'd115; b = 8'd176;  #10 
a = 8'd115; b = 8'd177;  #10 
a = 8'd115; b = 8'd178;  #10 
a = 8'd115; b = 8'd179;  #10 
a = 8'd115; b = 8'd180;  #10 
a = 8'd115; b = 8'd181;  #10 
a = 8'd115; b = 8'd182;  #10 
a = 8'd115; b = 8'd183;  #10 
a = 8'd115; b = 8'd184;  #10 
a = 8'd115; b = 8'd185;  #10 
a = 8'd115; b = 8'd186;  #10 
a = 8'd115; b = 8'd187;  #10 
a = 8'd115; b = 8'd188;  #10 
a = 8'd115; b = 8'd189;  #10 
a = 8'd115; b = 8'd190;  #10 
a = 8'd115; b = 8'd191;  #10 
a = 8'd115; b = 8'd192;  #10 
a = 8'd115; b = 8'd193;  #10 
a = 8'd115; b = 8'd194;  #10 
a = 8'd115; b = 8'd195;  #10 
a = 8'd115; b = 8'd196;  #10 
a = 8'd115; b = 8'd197;  #10 
a = 8'd115; b = 8'd198;  #10 
a = 8'd115; b = 8'd199;  #10 
a = 8'd115; b = 8'd200;  #10 
a = 8'd115; b = 8'd201;  #10 
a = 8'd115; b = 8'd202;  #10 
a = 8'd115; b = 8'd203;  #10 
a = 8'd115; b = 8'd204;  #10 
a = 8'd115; b = 8'd205;  #10 
a = 8'd115; b = 8'd206;  #10 
a = 8'd115; b = 8'd207;  #10 
a = 8'd115; b = 8'd208;  #10 
a = 8'd115; b = 8'd209;  #10 
a = 8'd115; b = 8'd210;  #10 
a = 8'd115; b = 8'd211;  #10 
a = 8'd115; b = 8'd212;  #10 
a = 8'd115; b = 8'd213;  #10 
a = 8'd115; b = 8'd214;  #10 
a = 8'd115; b = 8'd215;  #10 
a = 8'd115; b = 8'd216;  #10 
a = 8'd115; b = 8'd217;  #10 
a = 8'd115; b = 8'd218;  #10 
a = 8'd115; b = 8'd219;  #10 
a = 8'd115; b = 8'd220;  #10 
a = 8'd115; b = 8'd221;  #10 
a = 8'd115; b = 8'd222;  #10 
a = 8'd115; b = 8'd223;  #10 
a = 8'd115; b = 8'd224;  #10 
a = 8'd115; b = 8'd225;  #10 
a = 8'd115; b = 8'd226;  #10 
a = 8'd115; b = 8'd227;  #10 
a = 8'd115; b = 8'd228;  #10 
a = 8'd115; b = 8'd229;  #10 
a = 8'd115; b = 8'd230;  #10 
a = 8'd115; b = 8'd231;  #10 
a = 8'd115; b = 8'd232;  #10 
a = 8'd115; b = 8'd233;  #10 
a = 8'd115; b = 8'd234;  #10 
a = 8'd115; b = 8'd235;  #10 
a = 8'd115; b = 8'd236;  #10 
a = 8'd115; b = 8'd237;  #10 
a = 8'd115; b = 8'd238;  #10 
a = 8'd115; b = 8'd239;  #10 
a = 8'd115; b = 8'd240;  #10 
a = 8'd115; b = 8'd241;  #10 
a = 8'd115; b = 8'd242;  #10 
a = 8'd115; b = 8'd243;  #10 
a = 8'd115; b = 8'd244;  #10 
a = 8'd115; b = 8'd245;  #10 
a = 8'd115; b = 8'd246;  #10 
a = 8'd115; b = 8'd247;  #10 
a = 8'd115; b = 8'd248;  #10 
a = 8'd115; b = 8'd249;  #10 
a = 8'd115; b = 8'd250;  #10 
a = 8'd115; b = 8'd251;  #10 
a = 8'd115; b = 8'd252;  #10 
a = 8'd115; b = 8'd253;  #10 
a = 8'd115; b = 8'd254;  #10 
a = 8'd115; b = 8'd255;  #10 
a = 8'd116; b = 8'd0;  #10 
a = 8'd116; b = 8'd1;  #10 
a = 8'd116; b = 8'd2;  #10 
a = 8'd116; b = 8'd3;  #10 
a = 8'd116; b = 8'd4;  #10 
a = 8'd116; b = 8'd5;  #10 
a = 8'd116; b = 8'd6;  #10 
a = 8'd116; b = 8'd7;  #10 
a = 8'd116; b = 8'd8;  #10 
a = 8'd116; b = 8'd9;  #10 
a = 8'd116; b = 8'd10;  #10 
a = 8'd116; b = 8'd11;  #10 
a = 8'd116; b = 8'd12;  #10 
a = 8'd116; b = 8'd13;  #10 
a = 8'd116; b = 8'd14;  #10 
a = 8'd116; b = 8'd15;  #10 
a = 8'd116; b = 8'd16;  #10 
a = 8'd116; b = 8'd17;  #10 
a = 8'd116; b = 8'd18;  #10 
a = 8'd116; b = 8'd19;  #10 
a = 8'd116; b = 8'd20;  #10 
a = 8'd116; b = 8'd21;  #10 
a = 8'd116; b = 8'd22;  #10 
a = 8'd116; b = 8'd23;  #10 
a = 8'd116; b = 8'd24;  #10 
a = 8'd116; b = 8'd25;  #10 
a = 8'd116; b = 8'd26;  #10 
a = 8'd116; b = 8'd27;  #10 
a = 8'd116; b = 8'd28;  #10 
a = 8'd116; b = 8'd29;  #10 
a = 8'd116; b = 8'd30;  #10 
a = 8'd116; b = 8'd31;  #10 
a = 8'd116; b = 8'd32;  #10 
a = 8'd116; b = 8'd33;  #10 
a = 8'd116; b = 8'd34;  #10 
a = 8'd116; b = 8'd35;  #10 
a = 8'd116; b = 8'd36;  #10 
a = 8'd116; b = 8'd37;  #10 
a = 8'd116; b = 8'd38;  #10 
a = 8'd116; b = 8'd39;  #10 
a = 8'd116; b = 8'd40;  #10 
a = 8'd116; b = 8'd41;  #10 
a = 8'd116; b = 8'd42;  #10 
a = 8'd116; b = 8'd43;  #10 
a = 8'd116; b = 8'd44;  #10 
a = 8'd116; b = 8'd45;  #10 
a = 8'd116; b = 8'd46;  #10 
a = 8'd116; b = 8'd47;  #10 
a = 8'd116; b = 8'd48;  #10 
a = 8'd116; b = 8'd49;  #10 
a = 8'd116; b = 8'd50;  #10 
a = 8'd116; b = 8'd51;  #10 
a = 8'd116; b = 8'd52;  #10 
a = 8'd116; b = 8'd53;  #10 
a = 8'd116; b = 8'd54;  #10 
a = 8'd116; b = 8'd55;  #10 
a = 8'd116; b = 8'd56;  #10 
a = 8'd116; b = 8'd57;  #10 
a = 8'd116; b = 8'd58;  #10 
a = 8'd116; b = 8'd59;  #10 
a = 8'd116; b = 8'd60;  #10 
a = 8'd116; b = 8'd61;  #10 
a = 8'd116; b = 8'd62;  #10 
a = 8'd116; b = 8'd63;  #10 
a = 8'd116; b = 8'd64;  #10 
a = 8'd116; b = 8'd65;  #10 
a = 8'd116; b = 8'd66;  #10 
a = 8'd116; b = 8'd67;  #10 
a = 8'd116; b = 8'd68;  #10 
a = 8'd116; b = 8'd69;  #10 
a = 8'd116; b = 8'd70;  #10 
a = 8'd116; b = 8'd71;  #10 
a = 8'd116; b = 8'd72;  #10 
a = 8'd116; b = 8'd73;  #10 
a = 8'd116; b = 8'd74;  #10 
a = 8'd116; b = 8'd75;  #10 
a = 8'd116; b = 8'd76;  #10 
a = 8'd116; b = 8'd77;  #10 
a = 8'd116; b = 8'd78;  #10 
a = 8'd116; b = 8'd79;  #10 
a = 8'd116; b = 8'd80;  #10 
a = 8'd116; b = 8'd81;  #10 
a = 8'd116; b = 8'd82;  #10 
a = 8'd116; b = 8'd83;  #10 
a = 8'd116; b = 8'd84;  #10 
a = 8'd116; b = 8'd85;  #10 
a = 8'd116; b = 8'd86;  #10 
a = 8'd116; b = 8'd87;  #10 
a = 8'd116; b = 8'd88;  #10 
a = 8'd116; b = 8'd89;  #10 
a = 8'd116; b = 8'd90;  #10 
a = 8'd116; b = 8'd91;  #10 
a = 8'd116; b = 8'd92;  #10 
a = 8'd116; b = 8'd93;  #10 
a = 8'd116; b = 8'd94;  #10 
a = 8'd116; b = 8'd95;  #10 
a = 8'd116; b = 8'd96;  #10 
a = 8'd116; b = 8'd97;  #10 
a = 8'd116; b = 8'd98;  #10 
a = 8'd116; b = 8'd99;  #10 
a = 8'd116; b = 8'd100;  #10 
a = 8'd116; b = 8'd101;  #10 
a = 8'd116; b = 8'd102;  #10 
a = 8'd116; b = 8'd103;  #10 
a = 8'd116; b = 8'd104;  #10 
a = 8'd116; b = 8'd105;  #10 
a = 8'd116; b = 8'd106;  #10 
a = 8'd116; b = 8'd107;  #10 
a = 8'd116; b = 8'd108;  #10 
a = 8'd116; b = 8'd109;  #10 
a = 8'd116; b = 8'd110;  #10 
a = 8'd116; b = 8'd111;  #10 
a = 8'd116; b = 8'd112;  #10 
a = 8'd116; b = 8'd113;  #10 
a = 8'd116; b = 8'd114;  #10 
a = 8'd116; b = 8'd115;  #10 
a = 8'd116; b = 8'd116;  #10 
a = 8'd116; b = 8'd117;  #10 
a = 8'd116; b = 8'd118;  #10 
a = 8'd116; b = 8'd119;  #10 
a = 8'd116; b = 8'd120;  #10 
a = 8'd116; b = 8'd121;  #10 
a = 8'd116; b = 8'd122;  #10 
a = 8'd116; b = 8'd123;  #10 
a = 8'd116; b = 8'd124;  #10 
a = 8'd116; b = 8'd125;  #10 
a = 8'd116; b = 8'd126;  #10 
a = 8'd116; b = 8'd127;  #10 
a = 8'd116; b = 8'd128;  #10 
a = 8'd116; b = 8'd129;  #10 
a = 8'd116; b = 8'd130;  #10 
a = 8'd116; b = 8'd131;  #10 
a = 8'd116; b = 8'd132;  #10 
a = 8'd116; b = 8'd133;  #10 
a = 8'd116; b = 8'd134;  #10 
a = 8'd116; b = 8'd135;  #10 
a = 8'd116; b = 8'd136;  #10 
a = 8'd116; b = 8'd137;  #10 
a = 8'd116; b = 8'd138;  #10 
a = 8'd116; b = 8'd139;  #10 
a = 8'd116; b = 8'd140;  #10 
a = 8'd116; b = 8'd141;  #10 
a = 8'd116; b = 8'd142;  #10 
a = 8'd116; b = 8'd143;  #10 
a = 8'd116; b = 8'd144;  #10 
a = 8'd116; b = 8'd145;  #10 
a = 8'd116; b = 8'd146;  #10 
a = 8'd116; b = 8'd147;  #10 
a = 8'd116; b = 8'd148;  #10 
a = 8'd116; b = 8'd149;  #10 
a = 8'd116; b = 8'd150;  #10 
a = 8'd116; b = 8'd151;  #10 
a = 8'd116; b = 8'd152;  #10 
a = 8'd116; b = 8'd153;  #10 
a = 8'd116; b = 8'd154;  #10 
a = 8'd116; b = 8'd155;  #10 
a = 8'd116; b = 8'd156;  #10 
a = 8'd116; b = 8'd157;  #10 
a = 8'd116; b = 8'd158;  #10 
a = 8'd116; b = 8'd159;  #10 
a = 8'd116; b = 8'd160;  #10 
a = 8'd116; b = 8'd161;  #10 
a = 8'd116; b = 8'd162;  #10 
a = 8'd116; b = 8'd163;  #10 
a = 8'd116; b = 8'd164;  #10 
a = 8'd116; b = 8'd165;  #10 
a = 8'd116; b = 8'd166;  #10 
a = 8'd116; b = 8'd167;  #10 
a = 8'd116; b = 8'd168;  #10 
a = 8'd116; b = 8'd169;  #10 
a = 8'd116; b = 8'd170;  #10 
a = 8'd116; b = 8'd171;  #10 
a = 8'd116; b = 8'd172;  #10 
a = 8'd116; b = 8'd173;  #10 
a = 8'd116; b = 8'd174;  #10 
a = 8'd116; b = 8'd175;  #10 
a = 8'd116; b = 8'd176;  #10 
a = 8'd116; b = 8'd177;  #10 
a = 8'd116; b = 8'd178;  #10 
a = 8'd116; b = 8'd179;  #10 
a = 8'd116; b = 8'd180;  #10 
a = 8'd116; b = 8'd181;  #10 
a = 8'd116; b = 8'd182;  #10 
a = 8'd116; b = 8'd183;  #10 
a = 8'd116; b = 8'd184;  #10 
a = 8'd116; b = 8'd185;  #10 
a = 8'd116; b = 8'd186;  #10 
a = 8'd116; b = 8'd187;  #10 
a = 8'd116; b = 8'd188;  #10 
a = 8'd116; b = 8'd189;  #10 
a = 8'd116; b = 8'd190;  #10 
a = 8'd116; b = 8'd191;  #10 
a = 8'd116; b = 8'd192;  #10 
a = 8'd116; b = 8'd193;  #10 
a = 8'd116; b = 8'd194;  #10 
a = 8'd116; b = 8'd195;  #10 
a = 8'd116; b = 8'd196;  #10 
a = 8'd116; b = 8'd197;  #10 
a = 8'd116; b = 8'd198;  #10 
a = 8'd116; b = 8'd199;  #10 
a = 8'd116; b = 8'd200;  #10 
a = 8'd116; b = 8'd201;  #10 
a = 8'd116; b = 8'd202;  #10 
a = 8'd116; b = 8'd203;  #10 
a = 8'd116; b = 8'd204;  #10 
a = 8'd116; b = 8'd205;  #10 
a = 8'd116; b = 8'd206;  #10 
a = 8'd116; b = 8'd207;  #10 
a = 8'd116; b = 8'd208;  #10 
a = 8'd116; b = 8'd209;  #10 
a = 8'd116; b = 8'd210;  #10 
a = 8'd116; b = 8'd211;  #10 
a = 8'd116; b = 8'd212;  #10 
a = 8'd116; b = 8'd213;  #10 
a = 8'd116; b = 8'd214;  #10 
a = 8'd116; b = 8'd215;  #10 
a = 8'd116; b = 8'd216;  #10 
a = 8'd116; b = 8'd217;  #10 
a = 8'd116; b = 8'd218;  #10 
a = 8'd116; b = 8'd219;  #10 
a = 8'd116; b = 8'd220;  #10 
a = 8'd116; b = 8'd221;  #10 
a = 8'd116; b = 8'd222;  #10 
a = 8'd116; b = 8'd223;  #10 
a = 8'd116; b = 8'd224;  #10 
a = 8'd116; b = 8'd225;  #10 
a = 8'd116; b = 8'd226;  #10 
a = 8'd116; b = 8'd227;  #10 
a = 8'd116; b = 8'd228;  #10 
a = 8'd116; b = 8'd229;  #10 
a = 8'd116; b = 8'd230;  #10 
a = 8'd116; b = 8'd231;  #10 
a = 8'd116; b = 8'd232;  #10 
a = 8'd116; b = 8'd233;  #10 
a = 8'd116; b = 8'd234;  #10 
a = 8'd116; b = 8'd235;  #10 
a = 8'd116; b = 8'd236;  #10 
a = 8'd116; b = 8'd237;  #10 
a = 8'd116; b = 8'd238;  #10 
a = 8'd116; b = 8'd239;  #10 
a = 8'd116; b = 8'd240;  #10 
a = 8'd116; b = 8'd241;  #10 
a = 8'd116; b = 8'd242;  #10 
a = 8'd116; b = 8'd243;  #10 
a = 8'd116; b = 8'd244;  #10 
a = 8'd116; b = 8'd245;  #10 
a = 8'd116; b = 8'd246;  #10 
a = 8'd116; b = 8'd247;  #10 
a = 8'd116; b = 8'd248;  #10 
a = 8'd116; b = 8'd249;  #10 
a = 8'd116; b = 8'd250;  #10 
a = 8'd116; b = 8'd251;  #10 
a = 8'd116; b = 8'd252;  #10 
a = 8'd116; b = 8'd253;  #10 
a = 8'd116; b = 8'd254;  #10 
a = 8'd116; b = 8'd255;  #10 
a = 8'd117; b = 8'd0;  #10 
a = 8'd117; b = 8'd1;  #10 
a = 8'd117; b = 8'd2;  #10 
a = 8'd117; b = 8'd3;  #10 
a = 8'd117; b = 8'd4;  #10 
a = 8'd117; b = 8'd5;  #10 
a = 8'd117; b = 8'd6;  #10 
a = 8'd117; b = 8'd7;  #10 
a = 8'd117; b = 8'd8;  #10 
a = 8'd117; b = 8'd9;  #10 
a = 8'd117; b = 8'd10;  #10 
a = 8'd117; b = 8'd11;  #10 
a = 8'd117; b = 8'd12;  #10 
a = 8'd117; b = 8'd13;  #10 
a = 8'd117; b = 8'd14;  #10 
a = 8'd117; b = 8'd15;  #10 
a = 8'd117; b = 8'd16;  #10 
a = 8'd117; b = 8'd17;  #10 
a = 8'd117; b = 8'd18;  #10 
a = 8'd117; b = 8'd19;  #10 
a = 8'd117; b = 8'd20;  #10 
a = 8'd117; b = 8'd21;  #10 
a = 8'd117; b = 8'd22;  #10 
a = 8'd117; b = 8'd23;  #10 
a = 8'd117; b = 8'd24;  #10 
a = 8'd117; b = 8'd25;  #10 
a = 8'd117; b = 8'd26;  #10 
a = 8'd117; b = 8'd27;  #10 
a = 8'd117; b = 8'd28;  #10 
a = 8'd117; b = 8'd29;  #10 
a = 8'd117; b = 8'd30;  #10 
a = 8'd117; b = 8'd31;  #10 
a = 8'd117; b = 8'd32;  #10 
a = 8'd117; b = 8'd33;  #10 
a = 8'd117; b = 8'd34;  #10 
a = 8'd117; b = 8'd35;  #10 
a = 8'd117; b = 8'd36;  #10 
a = 8'd117; b = 8'd37;  #10 
a = 8'd117; b = 8'd38;  #10 
a = 8'd117; b = 8'd39;  #10 
a = 8'd117; b = 8'd40;  #10 
a = 8'd117; b = 8'd41;  #10 
a = 8'd117; b = 8'd42;  #10 
a = 8'd117; b = 8'd43;  #10 
a = 8'd117; b = 8'd44;  #10 
a = 8'd117; b = 8'd45;  #10 
a = 8'd117; b = 8'd46;  #10 
a = 8'd117; b = 8'd47;  #10 
a = 8'd117; b = 8'd48;  #10 
a = 8'd117; b = 8'd49;  #10 
a = 8'd117; b = 8'd50;  #10 
a = 8'd117; b = 8'd51;  #10 
a = 8'd117; b = 8'd52;  #10 
a = 8'd117; b = 8'd53;  #10 
a = 8'd117; b = 8'd54;  #10 
a = 8'd117; b = 8'd55;  #10 
a = 8'd117; b = 8'd56;  #10 
a = 8'd117; b = 8'd57;  #10 
a = 8'd117; b = 8'd58;  #10 
a = 8'd117; b = 8'd59;  #10 
a = 8'd117; b = 8'd60;  #10 
a = 8'd117; b = 8'd61;  #10 
a = 8'd117; b = 8'd62;  #10 
a = 8'd117; b = 8'd63;  #10 
a = 8'd117; b = 8'd64;  #10 
a = 8'd117; b = 8'd65;  #10 
a = 8'd117; b = 8'd66;  #10 
a = 8'd117; b = 8'd67;  #10 
a = 8'd117; b = 8'd68;  #10 
a = 8'd117; b = 8'd69;  #10 
a = 8'd117; b = 8'd70;  #10 
a = 8'd117; b = 8'd71;  #10 
a = 8'd117; b = 8'd72;  #10 
a = 8'd117; b = 8'd73;  #10 
a = 8'd117; b = 8'd74;  #10 
a = 8'd117; b = 8'd75;  #10 
a = 8'd117; b = 8'd76;  #10 
a = 8'd117; b = 8'd77;  #10 
a = 8'd117; b = 8'd78;  #10 
a = 8'd117; b = 8'd79;  #10 
a = 8'd117; b = 8'd80;  #10 
a = 8'd117; b = 8'd81;  #10 
a = 8'd117; b = 8'd82;  #10 
a = 8'd117; b = 8'd83;  #10 
a = 8'd117; b = 8'd84;  #10 
a = 8'd117; b = 8'd85;  #10 
a = 8'd117; b = 8'd86;  #10 
a = 8'd117; b = 8'd87;  #10 
a = 8'd117; b = 8'd88;  #10 
a = 8'd117; b = 8'd89;  #10 
a = 8'd117; b = 8'd90;  #10 
a = 8'd117; b = 8'd91;  #10 
a = 8'd117; b = 8'd92;  #10 
a = 8'd117; b = 8'd93;  #10 
a = 8'd117; b = 8'd94;  #10 
a = 8'd117; b = 8'd95;  #10 
a = 8'd117; b = 8'd96;  #10 
a = 8'd117; b = 8'd97;  #10 
a = 8'd117; b = 8'd98;  #10 
a = 8'd117; b = 8'd99;  #10 
a = 8'd117; b = 8'd100;  #10 
a = 8'd117; b = 8'd101;  #10 
a = 8'd117; b = 8'd102;  #10 
a = 8'd117; b = 8'd103;  #10 
a = 8'd117; b = 8'd104;  #10 
a = 8'd117; b = 8'd105;  #10 
a = 8'd117; b = 8'd106;  #10 
a = 8'd117; b = 8'd107;  #10 
a = 8'd117; b = 8'd108;  #10 
a = 8'd117; b = 8'd109;  #10 
a = 8'd117; b = 8'd110;  #10 
a = 8'd117; b = 8'd111;  #10 
a = 8'd117; b = 8'd112;  #10 
a = 8'd117; b = 8'd113;  #10 
a = 8'd117; b = 8'd114;  #10 
a = 8'd117; b = 8'd115;  #10 
a = 8'd117; b = 8'd116;  #10 
a = 8'd117; b = 8'd117;  #10 
a = 8'd117; b = 8'd118;  #10 
a = 8'd117; b = 8'd119;  #10 
a = 8'd117; b = 8'd120;  #10 
a = 8'd117; b = 8'd121;  #10 
a = 8'd117; b = 8'd122;  #10 
a = 8'd117; b = 8'd123;  #10 
a = 8'd117; b = 8'd124;  #10 
a = 8'd117; b = 8'd125;  #10 
a = 8'd117; b = 8'd126;  #10 
a = 8'd117; b = 8'd127;  #10 
a = 8'd117; b = 8'd128;  #10 
a = 8'd117; b = 8'd129;  #10 
a = 8'd117; b = 8'd130;  #10 
a = 8'd117; b = 8'd131;  #10 
a = 8'd117; b = 8'd132;  #10 
a = 8'd117; b = 8'd133;  #10 
a = 8'd117; b = 8'd134;  #10 
a = 8'd117; b = 8'd135;  #10 
a = 8'd117; b = 8'd136;  #10 
a = 8'd117; b = 8'd137;  #10 
a = 8'd117; b = 8'd138;  #10 
a = 8'd117; b = 8'd139;  #10 
a = 8'd117; b = 8'd140;  #10 
a = 8'd117; b = 8'd141;  #10 
a = 8'd117; b = 8'd142;  #10 
a = 8'd117; b = 8'd143;  #10 
a = 8'd117; b = 8'd144;  #10 
a = 8'd117; b = 8'd145;  #10 
a = 8'd117; b = 8'd146;  #10 
a = 8'd117; b = 8'd147;  #10 
a = 8'd117; b = 8'd148;  #10 
a = 8'd117; b = 8'd149;  #10 
a = 8'd117; b = 8'd150;  #10 
a = 8'd117; b = 8'd151;  #10 
a = 8'd117; b = 8'd152;  #10 
a = 8'd117; b = 8'd153;  #10 
a = 8'd117; b = 8'd154;  #10 
a = 8'd117; b = 8'd155;  #10 
a = 8'd117; b = 8'd156;  #10 
a = 8'd117; b = 8'd157;  #10 
a = 8'd117; b = 8'd158;  #10 
a = 8'd117; b = 8'd159;  #10 
a = 8'd117; b = 8'd160;  #10 
a = 8'd117; b = 8'd161;  #10 
a = 8'd117; b = 8'd162;  #10 
a = 8'd117; b = 8'd163;  #10 
a = 8'd117; b = 8'd164;  #10 
a = 8'd117; b = 8'd165;  #10 
a = 8'd117; b = 8'd166;  #10 
a = 8'd117; b = 8'd167;  #10 
a = 8'd117; b = 8'd168;  #10 
a = 8'd117; b = 8'd169;  #10 
a = 8'd117; b = 8'd170;  #10 
a = 8'd117; b = 8'd171;  #10 
a = 8'd117; b = 8'd172;  #10 
a = 8'd117; b = 8'd173;  #10 
a = 8'd117; b = 8'd174;  #10 
a = 8'd117; b = 8'd175;  #10 
a = 8'd117; b = 8'd176;  #10 
a = 8'd117; b = 8'd177;  #10 
a = 8'd117; b = 8'd178;  #10 
a = 8'd117; b = 8'd179;  #10 
a = 8'd117; b = 8'd180;  #10 
a = 8'd117; b = 8'd181;  #10 
a = 8'd117; b = 8'd182;  #10 
a = 8'd117; b = 8'd183;  #10 
a = 8'd117; b = 8'd184;  #10 
a = 8'd117; b = 8'd185;  #10 
a = 8'd117; b = 8'd186;  #10 
a = 8'd117; b = 8'd187;  #10 
a = 8'd117; b = 8'd188;  #10 
a = 8'd117; b = 8'd189;  #10 
a = 8'd117; b = 8'd190;  #10 
a = 8'd117; b = 8'd191;  #10 
a = 8'd117; b = 8'd192;  #10 
a = 8'd117; b = 8'd193;  #10 
a = 8'd117; b = 8'd194;  #10 
a = 8'd117; b = 8'd195;  #10 
a = 8'd117; b = 8'd196;  #10 
a = 8'd117; b = 8'd197;  #10 
a = 8'd117; b = 8'd198;  #10 
a = 8'd117; b = 8'd199;  #10 
a = 8'd117; b = 8'd200;  #10 
a = 8'd117; b = 8'd201;  #10 
a = 8'd117; b = 8'd202;  #10 
a = 8'd117; b = 8'd203;  #10 
a = 8'd117; b = 8'd204;  #10 
a = 8'd117; b = 8'd205;  #10 
a = 8'd117; b = 8'd206;  #10 
a = 8'd117; b = 8'd207;  #10 
a = 8'd117; b = 8'd208;  #10 
a = 8'd117; b = 8'd209;  #10 
a = 8'd117; b = 8'd210;  #10 
a = 8'd117; b = 8'd211;  #10 
a = 8'd117; b = 8'd212;  #10 
a = 8'd117; b = 8'd213;  #10 
a = 8'd117; b = 8'd214;  #10 
a = 8'd117; b = 8'd215;  #10 
a = 8'd117; b = 8'd216;  #10 
a = 8'd117; b = 8'd217;  #10 
a = 8'd117; b = 8'd218;  #10 
a = 8'd117; b = 8'd219;  #10 
a = 8'd117; b = 8'd220;  #10 
a = 8'd117; b = 8'd221;  #10 
a = 8'd117; b = 8'd222;  #10 
a = 8'd117; b = 8'd223;  #10 
a = 8'd117; b = 8'd224;  #10 
a = 8'd117; b = 8'd225;  #10 
a = 8'd117; b = 8'd226;  #10 
a = 8'd117; b = 8'd227;  #10 
a = 8'd117; b = 8'd228;  #10 
a = 8'd117; b = 8'd229;  #10 
a = 8'd117; b = 8'd230;  #10 
a = 8'd117; b = 8'd231;  #10 
a = 8'd117; b = 8'd232;  #10 
a = 8'd117; b = 8'd233;  #10 
a = 8'd117; b = 8'd234;  #10 
a = 8'd117; b = 8'd235;  #10 
a = 8'd117; b = 8'd236;  #10 
a = 8'd117; b = 8'd237;  #10 
a = 8'd117; b = 8'd238;  #10 
a = 8'd117; b = 8'd239;  #10 
a = 8'd117; b = 8'd240;  #10 
a = 8'd117; b = 8'd241;  #10 
a = 8'd117; b = 8'd242;  #10 
a = 8'd117; b = 8'd243;  #10 
a = 8'd117; b = 8'd244;  #10 
a = 8'd117; b = 8'd245;  #10 
a = 8'd117; b = 8'd246;  #10 
a = 8'd117; b = 8'd247;  #10 
a = 8'd117; b = 8'd248;  #10 
a = 8'd117; b = 8'd249;  #10 
a = 8'd117; b = 8'd250;  #10 
a = 8'd117; b = 8'd251;  #10 
a = 8'd117; b = 8'd252;  #10 
a = 8'd117; b = 8'd253;  #10 
a = 8'd117; b = 8'd254;  #10 
a = 8'd117; b = 8'd255;  #10 
a = 8'd118; b = 8'd0;  #10 
a = 8'd118; b = 8'd1;  #10 
a = 8'd118; b = 8'd2;  #10 
a = 8'd118; b = 8'd3;  #10 
a = 8'd118; b = 8'd4;  #10 
a = 8'd118; b = 8'd5;  #10 
a = 8'd118; b = 8'd6;  #10 
a = 8'd118; b = 8'd7;  #10 
a = 8'd118; b = 8'd8;  #10 
a = 8'd118; b = 8'd9;  #10 
a = 8'd118; b = 8'd10;  #10 
a = 8'd118; b = 8'd11;  #10 
a = 8'd118; b = 8'd12;  #10 
a = 8'd118; b = 8'd13;  #10 
a = 8'd118; b = 8'd14;  #10 
a = 8'd118; b = 8'd15;  #10 
a = 8'd118; b = 8'd16;  #10 
a = 8'd118; b = 8'd17;  #10 
a = 8'd118; b = 8'd18;  #10 
a = 8'd118; b = 8'd19;  #10 
a = 8'd118; b = 8'd20;  #10 
a = 8'd118; b = 8'd21;  #10 
a = 8'd118; b = 8'd22;  #10 
a = 8'd118; b = 8'd23;  #10 
a = 8'd118; b = 8'd24;  #10 
a = 8'd118; b = 8'd25;  #10 
a = 8'd118; b = 8'd26;  #10 
a = 8'd118; b = 8'd27;  #10 
a = 8'd118; b = 8'd28;  #10 
a = 8'd118; b = 8'd29;  #10 
a = 8'd118; b = 8'd30;  #10 
a = 8'd118; b = 8'd31;  #10 
a = 8'd118; b = 8'd32;  #10 
a = 8'd118; b = 8'd33;  #10 
a = 8'd118; b = 8'd34;  #10 
a = 8'd118; b = 8'd35;  #10 
a = 8'd118; b = 8'd36;  #10 
a = 8'd118; b = 8'd37;  #10 
a = 8'd118; b = 8'd38;  #10 
a = 8'd118; b = 8'd39;  #10 
a = 8'd118; b = 8'd40;  #10 
a = 8'd118; b = 8'd41;  #10 
a = 8'd118; b = 8'd42;  #10 
a = 8'd118; b = 8'd43;  #10 
a = 8'd118; b = 8'd44;  #10 
a = 8'd118; b = 8'd45;  #10 
a = 8'd118; b = 8'd46;  #10 
a = 8'd118; b = 8'd47;  #10 
a = 8'd118; b = 8'd48;  #10 
a = 8'd118; b = 8'd49;  #10 
a = 8'd118; b = 8'd50;  #10 
a = 8'd118; b = 8'd51;  #10 
a = 8'd118; b = 8'd52;  #10 
a = 8'd118; b = 8'd53;  #10 
a = 8'd118; b = 8'd54;  #10 
a = 8'd118; b = 8'd55;  #10 
a = 8'd118; b = 8'd56;  #10 
a = 8'd118; b = 8'd57;  #10 
a = 8'd118; b = 8'd58;  #10 
a = 8'd118; b = 8'd59;  #10 
a = 8'd118; b = 8'd60;  #10 
a = 8'd118; b = 8'd61;  #10 
a = 8'd118; b = 8'd62;  #10 
a = 8'd118; b = 8'd63;  #10 
a = 8'd118; b = 8'd64;  #10 
a = 8'd118; b = 8'd65;  #10 
a = 8'd118; b = 8'd66;  #10 
a = 8'd118; b = 8'd67;  #10 
a = 8'd118; b = 8'd68;  #10 
a = 8'd118; b = 8'd69;  #10 
a = 8'd118; b = 8'd70;  #10 
a = 8'd118; b = 8'd71;  #10 
a = 8'd118; b = 8'd72;  #10 
a = 8'd118; b = 8'd73;  #10 
a = 8'd118; b = 8'd74;  #10 
a = 8'd118; b = 8'd75;  #10 
a = 8'd118; b = 8'd76;  #10 
a = 8'd118; b = 8'd77;  #10 
a = 8'd118; b = 8'd78;  #10 
a = 8'd118; b = 8'd79;  #10 
a = 8'd118; b = 8'd80;  #10 
a = 8'd118; b = 8'd81;  #10 
a = 8'd118; b = 8'd82;  #10 
a = 8'd118; b = 8'd83;  #10 
a = 8'd118; b = 8'd84;  #10 
a = 8'd118; b = 8'd85;  #10 
a = 8'd118; b = 8'd86;  #10 
a = 8'd118; b = 8'd87;  #10 
a = 8'd118; b = 8'd88;  #10 
a = 8'd118; b = 8'd89;  #10 
a = 8'd118; b = 8'd90;  #10 
a = 8'd118; b = 8'd91;  #10 
a = 8'd118; b = 8'd92;  #10 
a = 8'd118; b = 8'd93;  #10 
a = 8'd118; b = 8'd94;  #10 
a = 8'd118; b = 8'd95;  #10 
a = 8'd118; b = 8'd96;  #10 
a = 8'd118; b = 8'd97;  #10 
a = 8'd118; b = 8'd98;  #10 
a = 8'd118; b = 8'd99;  #10 
a = 8'd118; b = 8'd100;  #10 
a = 8'd118; b = 8'd101;  #10 
a = 8'd118; b = 8'd102;  #10 
a = 8'd118; b = 8'd103;  #10 
a = 8'd118; b = 8'd104;  #10 
a = 8'd118; b = 8'd105;  #10 
a = 8'd118; b = 8'd106;  #10 
a = 8'd118; b = 8'd107;  #10 
a = 8'd118; b = 8'd108;  #10 
a = 8'd118; b = 8'd109;  #10 
a = 8'd118; b = 8'd110;  #10 
a = 8'd118; b = 8'd111;  #10 
a = 8'd118; b = 8'd112;  #10 
a = 8'd118; b = 8'd113;  #10 
a = 8'd118; b = 8'd114;  #10 
a = 8'd118; b = 8'd115;  #10 
a = 8'd118; b = 8'd116;  #10 
a = 8'd118; b = 8'd117;  #10 
a = 8'd118; b = 8'd118;  #10 
a = 8'd118; b = 8'd119;  #10 
a = 8'd118; b = 8'd120;  #10 
a = 8'd118; b = 8'd121;  #10 
a = 8'd118; b = 8'd122;  #10 
a = 8'd118; b = 8'd123;  #10 
a = 8'd118; b = 8'd124;  #10 
a = 8'd118; b = 8'd125;  #10 
a = 8'd118; b = 8'd126;  #10 
a = 8'd118; b = 8'd127;  #10 
a = 8'd118; b = 8'd128;  #10 
a = 8'd118; b = 8'd129;  #10 
a = 8'd118; b = 8'd130;  #10 
a = 8'd118; b = 8'd131;  #10 
a = 8'd118; b = 8'd132;  #10 
a = 8'd118; b = 8'd133;  #10 
a = 8'd118; b = 8'd134;  #10 
a = 8'd118; b = 8'd135;  #10 
a = 8'd118; b = 8'd136;  #10 
a = 8'd118; b = 8'd137;  #10 
a = 8'd118; b = 8'd138;  #10 
a = 8'd118; b = 8'd139;  #10 
a = 8'd118; b = 8'd140;  #10 
a = 8'd118; b = 8'd141;  #10 
a = 8'd118; b = 8'd142;  #10 
a = 8'd118; b = 8'd143;  #10 
a = 8'd118; b = 8'd144;  #10 
a = 8'd118; b = 8'd145;  #10 
a = 8'd118; b = 8'd146;  #10 
a = 8'd118; b = 8'd147;  #10 
a = 8'd118; b = 8'd148;  #10 
a = 8'd118; b = 8'd149;  #10 
a = 8'd118; b = 8'd150;  #10 
a = 8'd118; b = 8'd151;  #10 
a = 8'd118; b = 8'd152;  #10 
a = 8'd118; b = 8'd153;  #10 
a = 8'd118; b = 8'd154;  #10 
a = 8'd118; b = 8'd155;  #10 
a = 8'd118; b = 8'd156;  #10 
a = 8'd118; b = 8'd157;  #10 
a = 8'd118; b = 8'd158;  #10 
a = 8'd118; b = 8'd159;  #10 
a = 8'd118; b = 8'd160;  #10 
a = 8'd118; b = 8'd161;  #10 
a = 8'd118; b = 8'd162;  #10 
a = 8'd118; b = 8'd163;  #10 
a = 8'd118; b = 8'd164;  #10 
a = 8'd118; b = 8'd165;  #10 
a = 8'd118; b = 8'd166;  #10 
a = 8'd118; b = 8'd167;  #10 
a = 8'd118; b = 8'd168;  #10 
a = 8'd118; b = 8'd169;  #10 
a = 8'd118; b = 8'd170;  #10 
a = 8'd118; b = 8'd171;  #10 
a = 8'd118; b = 8'd172;  #10 
a = 8'd118; b = 8'd173;  #10 
a = 8'd118; b = 8'd174;  #10 
a = 8'd118; b = 8'd175;  #10 
a = 8'd118; b = 8'd176;  #10 
a = 8'd118; b = 8'd177;  #10 
a = 8'd118; b = 8'd178;  #10 
a = 8'd118; b = 8'd179;  #10 
a = 8'd118; b = 8'd180;  #10 
a = 8'd118; b = 8'd181;  #10 
a = 8'd118; b = 8'd182;  #10 
a = 8'd118; b = 8'd183;  #10 
a = 8'd118; b = 8'd184;  #10 
a = 8'd118; b = 8'd185;  #10 
a = 8'd118; b = 8'd186;  #10 
a = 8'd118; b = 8'd187;  #10 
a = 8'd118; b = 8'd188;  #10 
a = 8'd118; b = 8'd189;  #10 
a = 8'd118; b = 8'd190;  #10 
a = 8'd118; b = 8'd191;  #10 
a = 8'd118; b = 8'd192;  #10 
a = 8'd118; b = 8'd193;  #10 
a = 8'd118; b = 8'd194;  #10 
a = 8'd118; b = 8'd195;  #10 
a = 8'd118; b = 8'd196;  #10 
a = 8'd118; b = 8'd197;  #10 
a = 8'd118; b = 8'd198;  #10 
a = 8'd118; b = 8'd199;  #10 
a = 8'd118; b = 8'd200;  #10 
a = 8'd118; b = 8'd201;  #10 
a = 8'd118; b = 8'd202;  #10 
a = 8'd118; b = 8'd203;  #10 
a = 8'd118; b = 8'd204;  #10 
a = 8'd118; b = 8'd205;  #10 
a = 8'd118; b = 8'd206;  #10 
a = 8'd118; b = 8'd207;  #10 
a = 8'd118; b = 8'd208;  #10 
a = 8'd118; b = 8'd209;  #10 
a = 8'd118; b = 8'd210;  #10 
a = 8'd118; b = 8'd211;  #10 
a = 8'd118; b = 8'd212;  #10 
a = 8'd118; b = 8'd213;  #10 
a = 8'd118; b = 8'd214;  #10 
a = 8'd118; b = 8'd215;  #10 
a = 8'd118; b = 8'd216;  #10 
a = 8'd118; b = 8'd217;  #10 
a = 8'd118; b = 8'd218;  #10 
a = 8'd118; b = 8'd219;  #10 
a = 8'd118; b = 8'd220;  #10 
a = 8'd118; b = 8'd221;  #10 
a = 8'd118; b = 8'd222;  #10 
a = 8'd118; b = 8'd223;  #10 
a = 8'd118; b = 8'd224;  #10 
a = 8'd118; b = 8'd225;  #10 
a = 8'd118; b = 8'd226;  #10 
a = 8'd118; b = 8'd227;  #10 
a = 8'd118; b = 8'd228;  #10 
a = 8'd118; b = 8'd229;  #10 
a = 8'd118; b = 8'd230;  #10 
a = 8'd118; b = 8'd231;  #10 
a = 8'd118; b = 8'd232;  #10 
a = 8'd118; b = 8'd233;  #10 
a = 8'd118; b = 8'd234;  #10 
a = 8'd118; b = 8'd235;  #10 
a = 8'd118; b = 8'd236;  #10 
a = 8'd118; b = 8'd237;  #10 
a = 8'd118; b = 8'd238;  #10 
a = 8'd118; b = 8'd239;  #10 
a = 8'd118; b = 8'd240;  #10 
a = 8'd118; b = 8'd241;  #10 
a = 8'd118; b = 8'd242;  #10 
a = 8'd118; b = 8'd243;  #10 
a = 8'd118; b = 8'd244;  #10 
a = 8'd118; b = 8'd245;  #10 
a = 8'd118; b = 8'd246;  #10 
a = 8'd118; b = 8'd247;  #10 
a = 8'd118; b = 8'd248;  #10 
a = 8'd118; b = 8'd249;  #10 
a = 8'd118; b = 8'd250;  #10 
a = 8'd118; b = 8'd251;  #10 
a = 8'd118; b = 8'd252;  #10 
a = 8'd118; b = 8'd253;  #10 
a = 8'd118; b = 8'd254;  #10 
a = 8'd118; b = 8'd255;  #10 
a = 8'd119; b = 8'd0;  #10 
a = 8'd119; b = 8'd1;  #10 
a = 8'd119; b = 8'd2;  #10 
a = 8'd119; b = 8'd3;  #10 
a = 8'd119; b = 8'd4;  #10 
a = 8'd119; b = 8'd5;  #10 
a = 8'd119; b = 8'd6;  #10 
a = 8'd119; b = 8'd7;  #10 
a = 8'd119; b = 8'd8;  #10 
a = 8'd119; b = 8'd9;  #10 
a = 8'd119; b = 8'd10;  #10 
a = 8'd119; b = 8'd11;  #10 
a = 8'd119; b = 8'd12;  #10 
a = 8'd119; b = 8'd13;  #10 
a = 8'd119; b = 8'd14;  #10 
a = 8'd119; b = 8'd15;  #10 
a = 8'd119; b = 8'd16;  #10 
a = 8'd119; b = 8'd17;  #10 
a = 8'd119; b = 8'd18;  #10 
a = 8'd119; b = 8'd19;  #10 
a = 8'd119; b = 8'd20;  #10 
a = 8'd119; b = 8'd21;  #10 
a = 8'd119; b = 8'd22;  #10 
a = 8'd119; b = 8'd23;  #10 
a = 8'd119; b = 8'd24;  #10 
a = 8'd119; b = 8'd25;  #10 
a = 8'd119; b = 8'd26;  #10 
a = 8'd119; b = 8'd27;  #10 
a = 8'd119; b = 8'd28;  #10 
a = 8'd119; b = 8'd29;  #10 
a = 8'd119; b = 8'd30;  #10 
a = 8'd119; b = 8'd31;  #10 
a = 8'd119; b = 8'd32;  #10 
a = 8'd119; b = 8'd33;  #10 
a = 8'd119; b = 8'd34;  #10 
a = 8'd119; b = 8'd35;  #10 
a = 8'd119; b = 8'd36;  #10 
a = 8'd119; b = 8'd37;  #10 
a = 8'd119; b = 8'd38;  #10 
a = 8'd119; b = 8'd39;  #10 
a = 8'd119; b = 8'd40;  #10 
a = 8'd119; b = 8'd41;  #10 
a = 8'd119; b = 8'd42;  #10 
a = 8'd119; b = 8'd43;  #10 
a = 8'd119; b = 8'd44;  #10 
a = 8'd119; b = 8'd45;  #10 
a = 8'd119; b = 8'd46;  #10 
a = 8'd119; b = 8'd47;  #10 
a = 8'd119; b = 8'd48;  #10 
a = 8'd119; b = 8'd49;  #10 
a = 8'd119; b = 8'd50;  #10 
a = 8'd119; b = 8'd51;  #10 
a = 8'd119; b = 8'd52;  #10 
a = 8'd119; b = 8'd53;  #10 
a = 8'd119; b = 8'd54;  #10 
a = 8'd119; b = 8'd55;  #10 
a = 8'd119; b = 8'd56;  #10 
a = 8'd119; b = 8'd57;  #10 
a = 8'd119; b = 8'd58;  #10 
a = 8'd119; b = 8'd59;  #10 
a = 8'd119; b = 8'd60;  #10 
a = 8'd119; b = 8'd61;  #10 
a = 8'd119; b = 8'd62;  #10 
a = 8'd119; b = 8'd63;  #10 
a = 8'd119; b = 8'd64;  #10 
a = 8'd119; b = 8'd65;  #10 
a = 8'd119; b = 8'd66;  #10 
a = 8'd119; b = 8'd67;  #10 
a = 8'd119; b = 8'd68;  #10 
a = 8'd119; b = 8'd69;  #10 
a = 8'd119; b = 8'd70;  #10 
a = 8'd119; b = 8'd71;  #10 
a = 8'd119; b = 8'd72;  #10 
a = 8'd119; b = 8'd73;  #10 
a = 8'd119; b = 8'd74;  #10 
a = 8'd119; b = 8'd75;  #10 
a = 8'd119; b = 8'd76;  #10 
a = 8'd119; b = 8'd77;  #10 
a = 8'd119; b = 8'd78;  #10 
a = 8'd119; b = 8'd79;  #10 
a = 8'd119; b = 8'd80;  #10 
a = 8'd119; b = 8'd81;  #10 
a = 8'd119; b = 8'd82;  #10 
a = 8'd119; b = 8'd83;  #10 
a = 8'd119; b = 8'd84;  #10 
a = 8'd119; b = 8'd85;  #10 
a = 8'd119; b = 8'd86;  #10 
a = 8'd119; b = 8'd87;  #10 
a = 8'd119; b = 8'd88;  #10 
a = 8'd119; b = 8'd89;  #10 
a = 8'd119; b = 8'd90;  #10 
a = 8'd119; b = 8'd91;  #10 
a = 8'd119; b = 8'd92;  #10 
a = 8'd119; b = 8'd93;  #10 
a = 8'd119; b = 8'd94;  #10 
a = 8'd119; b = 8'd95;  #10 
a = 8'd119; b = 8'd96;  #10 
a = 8'd119; b = 8'd97;  #10 
a = 8'd119; b = 8'd98;  #10 
a = 8'd119; b = 8'd99;  #10 
a = 8'd119; b = 8'd100;  #10 
a = 8'd119; b = 8'd101;  #10 
a = 8'd119; b = 8'd102;  #10 
a = 8'd119; b = 8'd103;  #10 
a = 8'd119; b = 8'd104;  #10 
a = 8'd119; b = 8'd105;  #10 
a = 8'd119; b = 8'd106;  #10 
a = 8'd119; b = 8'd107;  #10 
a = 8'd119; b = 8'd108;  #10 
a = 8'd119; b = 8'd109;  #10 
a = 8'd119; b = 8'd110;  #10 
a = 8'd119; b = 8'd111;  #10 
a = 8'd119; b = 8'd112;  #10 
a = 8'd119; b = 8'd113;  #10 
a = 8'd119; b = 8'd114;  #10 
a = 8'd119; b = 8'd115;  #10 
a = 8'd119; b = 8'd116;  #10 
a = 8'd119; b = 8'd117;  #10 
a = 8'd119; b = 8'd118;  #10 
a = 8'd119; b = 8'd119;  #10 
a = 8'd119; b = 8'd120;  #10 
a = 8'd119; b = 8'd121;  #10 
a = 8'd119; b = 8'd122;  #10 
a = 8'd119; b = 8'd123;  #10 
a = 8'd119; b = 8'd124;  #10 
a = 8'd119; b = 8'd125;  #10 
a = 8'd119; b = 8'd126;  #10 
a = 8'd119; b = 8'd127;  #10 
a = 8'd119; b = 8'd128;  #10 
a = 8'd119; b = 8'd129;  #10 
a = 8'd119; b = 8'd130;  #10 
a = 8'd119; b = 8'd131;  #10 
a = 8'd119; b = 8'd132;  #10 
a = 8'd119; b = 8'd133;  #10 
a = 8'd119; b = 8'd134;  #10 
a = 8'd119; b = 8'd135;  #10 
a = 8'd119; b = 8'd136;  #10 
a = 8'd119; b = 8'd137;  #10 
a = 8'd119; b = 8'd138;  #10 
a = 8'd119; b = 8'd139;  #10 
a = 8'd119; b = 8'd140;  #10 
a = 8'd119; b = 8'd141;  #10 
a = 8'd119; b = 8'd142;  #10 
a = 8'd119; b = 8'd143;  #10 
a = 8'd119; b = 8'd144;  #10 
a = 8'd119; b = 8'd145;  #10 
a = 8'd119; b = 8'd146;  #10 
a = 8'd119; b = 8'd147;  #10 
a = 8'd119; b = 8'd148;  #10 
a = 8'd119; b = 8'd149;  #10 
a = 8'd119; b = 8'd150;  #10 
a = 8'd119; b = 8'd151;  #10 
a = 8'd119; b = 8'd152;  #10 
a = 8'd119; b = 8'd153;  #10 
a = 8'd119; b = 8'd154;  #10 
a = 8'd119; b = 8'd155;  #10 
a = 8'd119; b = 8'd156;  #10 
a = 8'd119; b = 8'd157;  #10 
a = 8'd119; b = 8'd158;  #10 
a = 8'd119; b = 8'd159;  #10 
a = 8'd119; b = 8'd160;  #10 
a = 8'd119; b = 8'd161;  #10 
a = 8'd119; b = 8'd162;  #10 
a = 8'd119; b = 8'd163;  #10 
a = 8'd119; b = 8'd164;  #10 
a = 8'd119; b = 8'd165;  #10 
a = 8'd119; b = 8'd166;  #10 
a = 8'd119; b = 8'd167;  #10 
a = 8'd119; b = 8'd168;  #10 
a = 8'd119; b = 8'd169;  #10 
a = 8'd119; b = 8'd170;  #10 
a = 8'd119; b = 8'd171;  #10 
a = 8'd119; b = 8'd172;  #10 
a = 8'd119; b = 8'd173;  #10 
a = 8'd119; b = 8'd174;  #10 
a = 8'd119; b = 8'd175;  #10 
a = 8'd119; b = 8'd176;  #10 
a = 8'd119; b = 8'd177;  #10 
a = 8'd119; b = 8'd178;  #10 
a = 8'd119; b = 8'd179;  #10 
a = 8'd119; b = 8'd180;  #10 
a = 8'd119; b = 8'd181;  #10 
a = 8'd119; b = 8'd182;  #10 
a = 8'd119; b = 8'd183;  #10 
a = 8'd119; b = 8'd184;  #10 
a = 8'd119; b = 8'd185;  #10 
a = 8'd119; b = 8'd186;  #10 
a = 8'd119; b = 8'd187;  #10 
a = 8'd119; b = 8'd188;  #10 
a = 8'd119; b = 8'd189;  #10 
a = 8'd119; b = 8'd190;  #10 
a = 8'd119; b = 8'd191;  #10 
a = 8'd119; b = 8'd192;  #10 
a = 8'd119; b = 8'd193;  #10 
a = 8'd119; b = 8'd194;  #10 
a = 8'd119; b = 8'd195;  #10 
a = 8'd119; b = 8'd196;  #10 
a = 8'd119; b = 8'd197;  #10 
a = 8'd119; b = 8'd198;  #10 
a = 8'd119; b = 8'd199;  #10 
a = 8'd119; b = 8'd200;  #10 
a = 8'd119; b = 8'd201;  #10 
a = 8'd119; b = 8'd202;  #10 
a = 8'd119; b = 8'd203;  #10 
a = 8'd119; b = 8'd204;  #10 
a = 8'd119; b = 8'd205;  #10 
a = 8'd119; b = 8'd206;  #10 
a = 8'd119; b = 8'd207;  #10 
a = 8'd119; b = 8'd208;  #10 
a = 8'd119; b = 8'd209;  #10 
a = 8'd119; b = 8'd210;  #10 
a = 8'd119; b = 8'd211;  #10 
a = 8'd119; b = 8'd212;  #10 
a = 8'd119; b = 8'd213;  #10 
a = 8'd119; b = 8'd214;  #10 
a = 8'd119; b = 8'd215;  #10 
a = 8'd119; b = 8'd216;  #10 
a = 8'd119; b = 8'd217;  #10 
a = 8'd119; b = 8'd218;  #10 
a = 8'd119; b = 8'd219;  #10 
a = 8'd119; b = 8'd220;  #10 
a = 8'd119; b = 8'd221;  #10 
a = 8'd119; b = 8'd222;  #10 
a = 8'd119; b = 8'd223;  #10 
a = 8'd119; b = 8'd224;  #10 
a = 8'd119; b = 8'd225;  #10 
a = 8'd119; b = 8'd226;  #10 
a = 8'd119; b = 8'd227;  #10 
a = 8'd119; b = 8'd228;  #10 
a = 8'd119; b = 8'd229;  #10 
a = 8'd119; b = 8'd230;  #10 
a = 8'd119; b = 8'd231;  #10 
a = 8'd119; b = 8'd232;  #10 
a = 8'd119; b = 8'd233;  #10 
a = 8'd119; b = 8'd234;  #10 
a = 8'd119; b = 8'd235;  #10 
a = 8'd119; b = 8'd236;  #10 
a = 8'd119; b = 8'd237;  #10 
a = 8'd119; b = 8'd238;  #10 
a = 8'd119; b = 8'd239;  #10 
a = 8'd119; b = 8'd240;  #10 
a = 8'd119; b = 8'd241;  #10 
a = 8'd119; b = 8'd242;  #10 
a = 8'd119; b = 8'd243;  #10 
a = 8'd119; b = 8'd244;  #10 
a = 8'd119; b = 8'd245;  #10 
a = 8'd119; b = 8'd246;  #10 
a = 8'd119; b = 8'd247;  #10 
a = 8'd119; b = 8'd248;  #10 
a = 8'd119; b = 8'd249;  #10 
a = 8'd119; b = 8'd250;  #10 
a = 8'd119; b = 8'd251;  #10 
a = 8'd119; b = 8'd252;  #10 
a = 8'd119; b = 8'd253;  #10 
a = 8'd119; b = 8'd254;  #10 
a = 8'd119; b = 8'd255;  #10 
a = 8'd120; b = 8'd0;  #10 
a = 8'd120; b = 8'd1;  #10 
a = 8'd120; b = 8'd2;  #10 
a = 8'd120; b = 8'd3;  #10 
a = 8'd120; b = 8'd4;  #10 
a = 8'd120; b = 8'd5;  #10 
a = 8'd120; b = 8'd6;  #10 
a = 8'd120; b = 8'd7;  #10 
a = 8'd120; b = 8'd8;  #10 
a = 8'd120; b = 8'd9;  #10 
a = 8'd120; b = 8'd10;  #10 
a = 8'd120; b = 8'd11;  #10 
a = 8'd120; b = 8'd12;  #10 
a = 8'd120; b = 8'd13;  #10 
a = 8'd120; b = 8'd14;  #10 
a = 8'd120; b = 8'd15;  #10 
a = 8'd120; b = 8'd16;  #10 
a = 8'd120; b = 8'd17;  #10 
a = 8'd120; b = 8'd18;  #10 
a = 8'd120; b = 8'd19;  #10 
a = 8'd120; b = 8'd20;  #10 
a = 8'd120; b = 8'd21;  #10 
a = 8'd120; b = 8'd22;  #10 
a = 8'd120; b = 8'd23;  #10 
a = 8'd120; b = 8'd24;  #10 
a = 8'd120; b = 8'd25;  #10 
a = 8'd120; b = 8'd26;  #10 
a = 8'd120; b = 8'd27;  #10 
a = 8'd120; b = 8'd28;  #10 
a = 8'd120; b = 8'd29;  #10 
a = 8'd120; b = 8'd30;  #10 
a = 8'd120; b = 8'd31;  #10 
a = 8'd120; b = 8'd32;  #10 
a = 8'd120; b = 8'd33;  #10 
a = 8'd120; b = 8'd34;  #10 
a = 8'd120; b = 8'd35;  #10 
a = 8'd120; b = 8'd36;  #10 
a = 8'd120; b = 8'd37;  #10 
a = 8'd120; b = 8'd38;  #10 
a = 8'd120; b = 8'd39;  #10 
a = 8'd120; b = 8'd40;  #10 
a = 8'd120; b = 8'd41;  #10 
a = 8'd120; b = 8'd42;  #10 
a = 8'd120; b = 8'd43;  #10 
a = 8'd120; b = 8'd44;  #10 
a = 8'd120; b = 8'd45;  #10 
a = 8'd120; b = 8'd46;  #10 
a = 8'd120; b = 8'd47;  #10 
a = 8'd120; b = 8'd48;  #10 
a = 8'd120; b = 8'd49;  #10 
a = 8'd120; b = 8'd50;  #10 
a = 8'd120; b = 8'd51;  #10 
a = 8'd120; b = 8'd52;  #10 
a = 8'd120; b = 8'd53;  #10 
a = 8'd120; b = 8'd54;  #10 
a = 8'd120; b = 8'd55;  #10 
a = 8'd120; b = 8'd56;  #10 
a = 8'd120; b = 8'd57;  #10 
a = 8'd120; b = 8'd58;  #10 
a = 8'd120; b = 8'd59;  #10 
a = 8'd120; b = 8'd60;  #10 
a = 8'd120; b = 8'd61;  #10 
a = 8'd120; b = 8'd62;  #10 
a = 8'd120; b = 8'd63;  #10 
a = 8'd120; b = 8'd64;  #10 
a = 8'd120; b = 8'd65;  #10 
a = 8'd120; b = 8'd66;  #10 
a = 8'd120; b = 8'd67;  #10 
a = 8'd120; b = 8'd68;  #10 
a = 8'd120; b = 8'd69;  #10 
a = 8'd120; b = 8'd70;  #10 
a = 8'd120; b = 8'd71;  #10 
a = 8'd120; b = 8'd72;  #10 
a = 8'd120; b = 8'd73;  #10 
a = 8'd120; b = 8'd74;  #10 
a = 8'd120; b = 8'd75;  #10 
a = 8'd120; b = 8'd76;  #10 
a = 8'd120; b = 8'd77;  #10 
a = 8'd120; b = 8'd78;  #10 
a = 8'd120; b = 8'd79;  #10 
a = 8'd120; b = 8'd80;  #10 
a = 8'd120; b = 8'd81;  #10 
a = 8'd120; b = 8'd82;  #10 
a = 8'd120; b = 8'd83;  #10 
a = 8'd120; b = 8'd84;  #10 
a = 8'd120; b = 8'd85;  #10 
a = 8'd120; b = 8'd86;  #10 
a = 8'd120; b = 8'd87;  #10 
a = 8'd120; b = 8'd88;  #10 
a = 8'd120; b = 8'd89;  #10 
a = 8'd120; b = 8'd90;  #10 
a = 8'd120; b = 8'd91;  #10 
a = 8'd120; b = 8'd92;  #10 
a = 8'd120; b = 8'd93;  #10 
a = 8'd120; b = 8'd94;  #10 
a = 8'd120; b = 8'd95;  #10 
a = 8'd120; b = 8'd96;  #10 
a = 8'd120; b = 8'd97;  #10 
a = 8'd120; b = 8'd98;  #10 
a = 8'd120; b = 8'd99;  #10 
a = 8'd120; b = 8'd100;  #10 
a = 8'd120; b = 8'd101;  #10 
a = 8'd120; b = 8'd102;  #10 
a = 8'd120; b = 8'd103;  #10 
a = 8'd120; b = 8'd104;  #10 
a = 8'd120; b = 8'd105;  #10 
a = 8'd120; b = 8'd106;  #10 
a = 8'd120; b = 8'd107;  #10 
a = 8'd120; b = 8'd108;  #10 
a = 8'd120; b = 8'd109;  #10 
a = 8'd120; b = 8'd110;  #10 
a = 8'd120; b = 8'd111;  #10 
a = 8'd120; b = 8'd112;  #10 
a = 8'd120; b = 8'd113;  #10 
a = 8'd120; b = 8'd114;  #10 
a = 8'd120; b = 8'd115;  #10 
a = 8'd120; b = 8'd116;  #10 
a = 8'd120; b = 8'd117;  #10 
a = 8'd120; b = 8'd118;  #10 
a = 8'd120; b = 8'd119;  #10 
a = 8'd120; b = 8'd120;  #10 
a = 8'd120; b = 8'd121;  #10 
a = 8'd120; b = 8'd122;  #10 
a = 8'd120; b = 8'd123;  #10 
a = 8'd120; b = 8'd124;  #10 
a = 8'd120; b = 8'd125;  #10 
a = 8'd120; b = 8'd126;  #10 
a = 8'd120; b = 8'd127;  #10 
a = 8'd120; b = 8'd128;  #10 
a = 8'd120; b = 8'd129;  #10 
a = 8'd120; b = 8'd130;  #10 
a = 8'd120; b = 8'd131;  #10 
a = 8'd120; b = 8'd132;  #10 
a = 8'd120; b = 8'd133;  #10 
a = 8'd120; b = 8'd134;  #10 
a = 8'd120; b = 8'd135;  #10 
a = 8'd120; b = 8'd136;  #10 
a = 8'd120; b = 8'd137;  #10 
a = 8'd120; b = 8'd138;  #10 
a = 8'd120; b = 8'd139;  #10 
a = 8'd120; b = 8'd140;  #10 
a = 8'd120; b = 8'd141;  #10 
a = 8'd120; b = 8'd142;  #10 
a = 8'd120; b = 8'd143;  #10 
a = 8'd120; b = 8'd144;  #10 
a = 8'd120; b = 8'd145;  #10 
a = 8'd120; b = 8'd146;  #10 
a = 8'd120; b = 8'd147;  #10 
a = 8'd120; b = 8'd148;  #10 
a = 8'd120; b = 8'd149;  #10 
a = 8'd120; b = 8'd150;  #10 
a = 8'd120; b = 8'd151;  #10 
a = 8'd120; b = 8'd152;  #10 
a = 8'd120; b = 8'd153;  #10 
a = 8'd120; b = 8'd154;  #10 
a = 8'd120; b = 8'd155;  #10 
a = 8'd120; b = 8'd156;  #10 
a = 8'd120; b = 8'd157;  #10 
a = 8'd120; b = 8'd158;  #10 
a = 8'd120; b = 8'd159;  #10 
a = 8'd120; b = 8'd160;  #10 
a = 8'd120; b = 8'd161;  #10 
a = 8'd120; b = 8'd162;  #10 
a = 8'd120; b = 8'd163;  #10 
a = 8'd120; b = 8'd164;  #10 
a = 8'd120; b = 8'd165;  #10 
a = 8'd120; b = 8'd166;  #10 
a = 8'd120; b = 8'd167;  #10 
a = 8'd120; b = 8'd168;  #10 
a = 8'd120; b = 8'd169;  #10 
a = 8'd120; b = 8'd170;  #10 
a = 8'd120; b = 8'd171;  #10 
a = 8'd120; b = 8'd172;  #10 
a = 8'd120; b = 8'd173;  #10 
a = 8'd120; b = 8'd174;  #10 
a = 8'd120; b = 8'd175;  #10 
a = 8'd120; b = 8'd176;  #10 
a = 8'd120; b = 8'd177;  #10 
a = 8'd120; b = 8'd178;  #10 
a = 8'd120; b = 8'd179;  #10 
a = 8'd120; b = 8'd180;  #10 
a = 8'd120; b = 8'd181;  #10 
a = 8'd120; b = 8'd182;  #10 
a = 8'd120; b = 8'd183;  #10 
a = 8'd120; b = 8'd184;  #10 
a = 8'd120; b = 8'd185;  #10 
a = 8'd120; b = 8'd186;  #10 
a = 8'd120; b = 8'd187;  #10 
a = 8'd120; b = 8'd188;  #10 
a = 8'd120; b = 8'd189;  #10 
a = 8'd120; b = 8'd190;  #10 
a = 8'd120; b = 8'd191;  #10 
a = 8'd120; b = 8'd192;  #10 
a = 8'd120; b = 8'd193;  #10 
a = 8'd120; b = 8'd194;  #10 
a = 8'd120; b = 8'd195;  #10 
a = 8'd120; b = 8'd196;  #10 
a = 8'd120; b = 8'd197;  #10 
a = 8'd120; b = 8'd198;  #10 
a = 8'd120; b = 8'd199;  #10 
a = 8'd120; b = 8'd200;  #10 
a = 8'd120; b = 8'd201;  #10 
a = 8'd120; b = 8'd202;  #10 
a = 8'd120; b = 8'd203;  #10 
a = 8'd120; b = 8'd204;  #10 
a = 8'd120; b = 8'd205;  #10 
a = 8'd120; b = 8'd206;  #10 
a = 8'd120; b = 8'd207;  #10 
a = 8'd120; b = 8'd208;  #10 
a = 8'd120; b = 8'd209;  #10 
a = 8'd120; b = 8'd210;  #10 
a = 8'd120; b = 8'd211;  #10 
a = 8'd120; b = 8'd212;  #10 
a = 8'd120; b = 8'd213;  #10 
a = 8'd120; b = 8'd214;  #10 
a = 8'd120; b = 8'd215;  #10 
a = 8'd120; b = 8'd216;  #10 
a = 8'd120; b = 8'd217;  #10 
a = 8'd120; b = 8'd218;  #10 
a = 8'd120; b = 8'd219;  #10 
a = 8'd120; b = 8'd220;  #10 
a = 8'd120; b = 8'd221;  #10 
a = 8'd120; b = 8'd222;  #10 
a = 8'd120; b = 8'd223;  #10 
a = 8'd120; b = 8'd224;  #10 
a = 8'd120; b = 8'd225;  #10 
a = 8'd120; b = 8'd226;  #10 
a = 8'd120; b = 8'd227;  #10 
a = 8'd120; b = 8'd228;  #10 
a = 8'd120; b = 8'd229;  #10 
a = 8'd120; b = 8'd230;  #10 
a = 8'd120; b = 8'd231;  #10 
a = 8'd120; b = 8'd232;  #10 
a = 8'd120; b = 8'd233;  #10 
a = 8'd120; b = 8'd234;  #10 
a = 8'd120; b = 8'd235;  #10 
a = 8'd120; b = 8'd236;  #10 
a = 8'd120; b = 8'd237;  #10 
a = 8'd120; b = 8'd238;  #10 
a = 8'd120; b = 8'd239;  #10 
a = 8'd120; b = 8'd240;  #10 
a = 8'd120; b = 8'd241;  #10 
a = 8'd120; b = 8'd242;  #10 
a = 8'd120; b = 8'd243;  #10 
a = 8'd120; b = 8'd244;  #10 
a = 8'd120; b = 8'd245;  #10 
a = 8'd120; b = 8'd246;  #10 
a = 8'd120; b = 8'd247;  #10 
a = 8'd120; b = 8'd248;  #10 
a = 8'd120; b = 8'd249;  #10 
a = 8'd120; b = 8'd250;  #10 
a = 8'd120; b = 8'd251;  #10 
a = 8'd120; b = 8'd252;  #10 
a = 8'd120; b = 8'd253;  #10 
a = 8'd120; b = 8'd254;  #10 
a = 8'd120; b = 8'd255;  #10 
a = 8'd121; b = 8'd0;  #10 
a = 8'd121; b = 8'd1;  #10 
a = 8'd121; b = 8'd2;  #10 
a = 8'd121; b = 8'd3;  #10 
a = 8'd121; b = 8'd4;  #10 
a = 8'd121; b = 8'd5;  #10 
a = 8'd121; b = 8'd6;  #10 
a = 8'd121; b = 8'd7;  #10 
a = 8'd121; b = 8'd8;  #10 
a = 8'd121; b = 8'd9;  #10 
a = 8'd121; b = 8'd10;  #10 
a = 8'd121; b = 8'd11;  #10 
a = 8'd121; b = 8'd12;  #10 
a = 8'd121; b = 8'd13;  #10 
a = 8'd121; b = 8'd14;  #10 
a = 8'd121; b = 8'd15;  #10 
a = 8'd121; b = 8'd16;  #10 
a = 8'd121; b = 8'd17;  #10 
a = 8'd121; b = 8'd18;  #10 
a = 8'd121; b = 8'd19;  #10 
a = 8'd121; b = 8'd20;  #10 
a = 8'd121; b = 8'd21;  #10 
a = 8'd121; b = 8'd22;  #10 
a = 8'd121; b = 8'd23;  #10 
a = 8'd121; b = 8'd24;  #10 
a = 8'd121; b = 8'd25;  #10 
a = 8'd121; b = 8'd26;  #10 
a = 8'd121; b = 8'd27;  #10 
a = 8'd121; b = 8'd28;  #10 
a = 8'd121; b = 8'd29;  #10 
a = 8'd121; b = 8'd30;  #10 
a = 8'd121; b = 8'd31;  #10 
a = 8'd121; b = 8'd32;  #10 
a = 8'd121; b = 8'd33;  #10 
a = 8'd121; b = 8'd34;  #10 
a = 8'd121; b = 8'd35;  #10 
a = 8'd121; b = 8'd36;  #10 
a = 8'd121; b = 8'd37;  #10 
a = 8'd121; b = 8'd38;  #10 
a = 8'd121; b = 8'd39;  #10 
a = 8'd121; b = 8'd40;  #10 
a = 8'd121; b = 8'd41;  #10 
a = 8'd121; b = 8'd42;  #10 
a = 8'd121; b = 8'd43;  #10 
a = 8'd121; b = 8'd44;  #10 
a = 8'd121; b = 8'd45;  #10 
a = 8'd121; b = 8'd46;  #10 
a = 8'd121; b = 8'd47;  #10 
a = 8'd121; b = 8'd48;  #10 
a = 8'd121; b = 8'd49;  #10 
a = 8'd121; b = 8'd50;  #10 
a = 8'd121; b = 8'd51;  #10 
a = 8'd121; b = 8'd52;  #10 
a = 8'd121; b = 8'd53;  #10 
a = 8'd121; b = 8'd54;  #10 
a = 8'd121; b = 8'd55;  #10 
a = 8'd121; b = 8'd56;  #10 
a = 8'd121; b = 8'd57;  #10 
a = 8'd121; b = 8'd58;  #10 
a = 8'd121; b = 8'd59;  #10 
a = 8'd121; b = 8'd60;  #10 
a = 8'd121; b = 8'd61;  #10 
a = 8'd121; b = 8'd62;  #10 
a = 8'd121; b = 8'd63;  #10 
a = 8'd121; b = 8'd64;  #10 
a = 8'd121; b = 8'd65;  #10 
a = 8'd121; b = 8'd66;  #10 
a = 8'd121; b = 8'd67;  #10 
a = 8'd121; b = 8'd68;  #10 
a = 8'd121; b = 8'd69;  #10 
a = 8'd121; b = 8'd70;  #10 
a = 8'd121; b = 8'd71;  #10 
a = 8'd121; b = 8'd72;  #10 
a = 8'd121; b = 8'd73;  #10 
a = 8'd121; b = 8'd74;  #10 
a = 8'd121; b = 8'd75;  #10 
a = 8'd121; b = 8'd76;  #10 
a = 8'd121; b = 8'd77;  #10 
a = 8'd121; b = 8'd78;  #10 
a = 8'd121; b = 8'd79;  #10 
a = 8'd121; b = 8'd80;  #10 
a = 8'd121; b = 8'd81;  #10 
a = 8'd121; b = 8'd82;  #10 
a = 8'd121; b = 8'd83;  #10 
a = 8'd121; b = 8'd84;  #10 
a = 8'd121; b = 8'd85;  #10 
a = 8'd121; b = 8'd86;  #10 
a = 8'd121; b = 8'd87;  #10 
a = 8'd121; b = 8'd88;  #10 
a = 8'd121; b = 8'd89;  #10 
a = 8'd121; b = 8'd90;  #10 
a = 8'd121; b = 8'd91;  #10 
a = 8'd121; b = 8'd92;  #10 
a = 8'd121; b = 8'd93;  #10 
a = 8'd121; b = 8'd94;  #10 
a = 8'd121; b = 8'd95;  #10 
a = 8'd121; b = 8'd96;  #10 
a = 8'd121; b = 8'd97;  #10 
a = 8'd121; b = 8'd98;  #10 
a = 8'd121; b = 8'd99;  #10 
a = 8'd121; b = 8'd100;  #10 
a = 8'd121; b = 8'd101;  #10 
a = 8'd121; b = 8'd102;  #10 
a = 8'd121; b = 8'd103;  #10 
a = 8'd121; b = 8'd104;  #10 
a = 8'd121; b = 8'd105;  #10 
a = 8'd121; b = 8'd106;  #10 
a = 8'd121; b = 8'd107;  #10 
a = 8'd121; b = 8'd108;  #10 
a = 8'd121; b = 8'd109;  #10 
a = 8'd121; b = 8'd110;  #10 
a = 8'd121; b = 8'd111;  #10 
a = 8'd121; b = 8'd112;  #10 
a = 8'd121; b = 8'd113;  #10 
a = 8'd121; b = 8'd114;  #10 
a = 8'd121; b = 8'd115;  #10 
a = 8'd121; b = 8'd116;  #10 
a = 8'd121; b = 8'd117;  #10 
a = 8'd121; b = 8'd118;  #10 
a = 8'd121; b = 8'd119;  #10 
a = 8'd121; b = 8'd120;  #10 
a = 8'd121; b = 8'd121;  #10 
a = 8'd121; b = 8'd122;  #10 
a = 8'd121; b = 8'd123;  #10 
a = 8'd121; b = 8'd124;  #10 
a = 8'd121; b = 8'd125;  #10 
a = 8'd121; b = 8'd126;  #10 
a = 8'd121; b = 8'd127;  #10 
a = 8'd121; b = 8'd128;  #10 
a = 8'd121; b = 8'd129;  #10 
a = 8'd121; b = 8'd130;  #10 
a = 8'd121; b = 8'd131;  #10 
a = 8'd121; b = 8'd132;  #10 
a = 8'd121; b = 8'd133;  #10 
a = 8'd121; b = 8'd134;  #10 
a = 8'd121; b = 8'd135;  #10 
a = 8'd121; b = 8'd136;  #10 
a = 8'd121; b = 8'd137;  #10 
a = 8'd121; b = 8'd138;  #10 
a = 8'd121; b = 8'd139;  #10 
a = 8'd121; b = 8'd140;  #10 
a = 8'd121; b = 8'd141;  #10 
a = 8'd121; b = 8'd142;  #10 
a = 8'd121; b = 8'd143;  #10 
a = 8'd121; b = 8'd144;  #10 
a = 8'd121; b = 8'd145;  #10 
a = 8'd121; b = 8'd146;  #10 
a = 8'd121; b = 8'd147;  #10 
a = 8'd121; b = 8'd148;  #10 
a = 8'd121; b = 8'd149;  #10 
a = 8'd121; b = 8'd150;  #10 
a = 8'd121; b = 8'd151;  #10 
a = 8'd121; b = 8'd152;  #10 
a = 8'd121; b = 8'd153;  #10 
a = 8'd121; b = 8'd154;  #10 
a = 8'd121; b = 8'd155;  #10 
a = 8'd121; b = 8'd156;  #10 
a = 8'd121; b = 8'd157;  #10 
a = 8'd121; b = 8'd158;  #10 
a = 8'd121; b = 8'd159;  #10 
a = 8'd121; b = 8'd160;  #10 
a = 8'd121; b = 8'd161;  #10 
a = 8'd121; b = 8'd162;  #10 
a = 8'd121; b = 8'd163;  #10 
a = 8'd121; b = 8'd164;  #10 
a = 8'd121; b = 8'd165;  #10 
a = 8'd121; b = 8'd166;  #10 
a = 8'd121; b = 8'd167;  #10 
a = 8'd121; b = 8'd168;  #10 
a = 8'd121; b = 8'd169;  #10 
a = 8'd121; b = 8'd170;  #10 
a = 8'd121; b = 8'd171;  #10 
a = 8'd121; b = 8'd172;  #10 
a = 8'd121; b = 8'd173;  #10 
a = 8'd121; b = 8'd174;  #10 
a = 8'd121; b = 8'd175;  #10 
a = 8'd121; b = 8'd176;  #10 
a = 8'd121; b = 8'd177;  #10 
a = 8'd121; b = 8'd178;  #10 
a = 8'd121; b = 8'd179;  #10 
a = 8'd121; b = 8'd180;  #10 
a = 8'd121; b = 8'd181;  #10 
a = 8'd121; b = 8'd182;  #10 
a = 8'd121; b = 8'd183;  #10 
a = 8'd121; b = 8'd184;  #10 
a = 8'd121; b = 8'd185;  #10 
a = 8'd121; b = 8'd186;  #10 
a = 8'd121; b = 8'd187;  #10 
a = 8'd121; b = 8'd188;  #10 
a = 8'd121; b = 8'd189;  #10 
a = 8'd121; b = 8'd190;  #10 
a = 8'd121; b = 8'd191;  #10 
a = 8'd121; b = 8'd192;  #10 
a = 8'd121; b = 8'd193;  #10 
a = 8'd121; b = 8'd194;  #10 
a = 8'd121; b = 8'd195;  #10 
a = 8'd121; b = 8'd196;  #10 
a = 8'd121; b = 8'd197;  #10 
a = 8'd121; b = 8'd198;  #10 
a = 8'd121; b = 8'd199;  #10 
a = 8'd121; b = 8'd200;  #10 
a = 8'd121; b = 8'd201;  #10 
a = 8'd121; b = 8'd202;  #10 
a = 8'd121; b = 8'd203;  #10 
a = 8'd121; b = 8'd204;  #10 
a = 8'd121; b = 8'd205;  #10 
a = 8'd121; b = 8'd206;  #10 
a = 8'd121; b = 8'd207;  #10 
a = 8'd121; b = 8'd208;  #10 
a = 8'd121; b = 8'd209;  #10 
a = 8'd121; b = 8'd210;  #10 
a = 8'd121; b = 8'd211;  #10 
a = 8'd121; b = 8'd212;  #10 
a = 8'd121; b = 8'd213;  #10 
a = 8'd121; b = 8'd214;  #10 
a = 8'd121; b = 8'd215;  #10 
a = 8'd121; b = 8'd216;  #10 
a = 8'd121; b = 8'd217;  #10 
a = 8'd121; b = 8'd218;  #10 
a = 8'd121; b = 8'd219;  #10 
a = 8'd121; b = 8'd220;  #10 
a = 8'd121; b = 8'd221;  #10 
a = 8'd121; b = 8'd222;  #10 
a = 8'd121; b = 8'd223;  #10 
a = 8'd121; b = 8'd224;  #10 
a = 8'd121; b = 8'd225;  #10 
a = 8'd121; b = 8'd226;  #10 
a = 8'd121; b = 8'd227;  #10 
a = 8'd121; b = 8'd228;  #10 
a = 8'd121; b = 8'd229;  #10 
a = 8'd121; b = 8'd230;  #10 
a = 8'd121; b = 8'd231;  #10 
a = 8'd121; b = 8'd232;  #10 
a = 8'd121; b = 8'd233;  #10 
a = 8'd121; b = 8'd234;  #10 
a = 8'd121; b = 8'd235;  #10 
a = 8'd121; b = 8'd236;  #10 
a = 8'd121; b = 8'd237;  #10 
a = 8'd121; b = 8'd238;  #10 
a = 8'd121; b = 8'd239;  #10 
a = 8'd121; b = 8'd240;  #10 
a = 8'd121; b = 8'd241;  #10 
a = 8'd121; b = 8'd242;  #10 
a = 8'd121; b = 8'd243;  #10 
a = 8'd121; b = 8'd244;  #10 
a = 8'd121; b = 8'd245;  #10 
a = 8'd121; b = 8'd246;  #10 
a = 8'd121; b = 8'd247;  #10 
a = 8'd121; b = 8'd248;  #10 
a = 8'd121; b = 8'd249;  #10 
a = 8'd121; b = 8'd250;  #10 
a = 8'd121; b = 8'd251;  #10 
a = 8'd121; b = 8'd252;  #10 
a = 8'd121; b = 8'd253;  #10 
a = 8'd121; b = 8'd254;  #10 
a = 8'd121; b = 8'd255;  #10 
a = 8'd122; b = 8'd0;  #10 
a = 8'd122; b = 8'd1;  #10 
a = 8'd122; b = 8'd2;  #10 
a = 8'd122; b = 8'd3;  #10 
a = 8'd122; b = 8'd4;  #10 
a = 8'd122; b = 8'd5;  #10 
a = 8'd122; b = 8'd6;  #10 
a = 8'd122; b = 8'd7;  #10 
a = 8'd122; b = 8'd8;  #10 
a = 8'd122; b = 8'd9;  #10 
a = 8'd122; b = 8'd10;  #10 
a = 8'd122; b = 8'd11;  #10 
a = 8'd122; b = 8'd12;  #10 
a = 8'd122; b = 8'd13;  #10 
a = 8'd122; b = 8'd14;  #10 
a = 8'd122; b = 8'd15;  #10 
a = 8'd122; b = 8'd16;  #10 
a = 8'd122; b = 8'd17;  #10 
a = 8'd122; b = 8'd18;  #10 
a = 8'd122; b = 8'd19;  #10 
a = 8'd122; b = 8'd20;  #10 
a = 8'd122; b = 8'd21;  #10 
a = 8'd122; b = 8'd22;  #10 
a = 8'd122; b = 8'd23;  #10 
a = 8'd122; b = 8'd24;  #10 
a = 8'd122; b = 8'd25;  #10 
a = 8'd122; b = 8'd26;  #10 
a = 8'd122; b = 8'd27;  #10 
a = 8'd122; b = 8'd28;  #10 
a = 8'd122; b = 8'd29;  #10 
a = 8'd122; b = 8'd30;  #10 
a = 8'd122; b = 8'd31;  #10 
a = 8'd122; b = 8'd32;  #10 
a = 8'd122; b = 8'd33;  #10 
a = 8'd122; b = 8'd34;  #10 
a = 8'd122; b = 8'd35;  #10 
a = 8'd122; b = 8'd36;  #10 
a = 8'd122; b = 8'd37;  #10 
a = 8'd122; b = 8'd38;  #10 
a = 8'd122; b = 8'd39;  #10 
a = 8'd122; b = 8'd40;  #10 
a = 8'd122; b = 8'd41;  #10 
a = 8'd122; b = 8'd42;  #10 
a = 8'd122; b = 8'd43;  #10 
a = 8'd122; b = 8'd44;  #10 
a = 8'd122; b = 8'd45;  #10 
a = 8'd122; b = 8'd46;  #10 
a = 8'd122; b = 8'd47;  #10 
a = 8'd122; b = 8'd48;  #10 
a = 8'd122; b = 8'd49;  #10 
a = 8'd122; b = 8'd50;  #10 
a = 8'd122; b = 8'd51;  #10 
a = 8'd122; b = 8'd52;  #10 
a = 8'd122; b = 8'd53;  #10 
a = 8'd122; b = 8'd54;  #10 
a = 8'd122; b = 8'd55;  #10 
a = 8'd122; b = 8'd56;  #10 
a = 8'd122; b = 8'd57;  #10 
a = 8'd122; b = 8'd58;  #10 
a = 8'd122; b = 8'd59;  #10 
a = 8'd122; b = 8'd60;  #10 
a = 8'd122; b = 8'd61;  #10 
a = 8'd122; b = 8'd62;  #10 
a = 8'd122; b = 8'd63;  #10 
a = 8'd122; b = 8'd64;  #10 
a = 8'd122; b = 8'd65;  #10 
a = 8'd122; b = 8'd66;  #10 
a = 8'd122; b = 8'd67;  #10 
a = 8'd122; b = 8'd68;  #10 
a = 8'd122; b = 8'd69;  #10 
a = 8'd122; b = 8'd70;  #10 
a = 8'd122; b = 8'd71;  #10 
a = 8'd122; b = 8'd72;  #10 
a = 8'd122; b = 8'd73;  #10 
a = 8'd122; b = 8'd74;  #10 
a = 8'd122; b = 8'd75;  #10 
a = 8'd122; b = 8'd76;  #10 
a = 8'd122; b = 8'd77;  #10 
a = 8'd122; b = 8'd78;  #10 
a = 8'd122; b = 8'd79;  #10 
a = 8'd122; b = 8'd80;  #10 
a = 8'd122; b = 8'd81;  #10 
a = 8'd122; b = 8'd82;  #10 
a = 8'd122; b = 8'd83;  #10 
a = 8'd122; b = 8'd84;  #10 
a = 8'd122; b = 8'd85;  #10 
a = 8'd122; b = 8'd86;  #10 
a = 8'd122; b = 8'd87;  #10 
a = 8'd122; b = 8'd88;  #10 
a = 8'd122; b = 8'd89;  #10 
a = 8'd122; b = 8'd90;  #10 
a = 8'd122; b = 8'd91;  #10 
a = 8'd122; b = 8'd92;  #10 
a = 8'd122; b = 8'd93;  #10 
a = 8'd122; b = 8'd94;  #10 
a = 8'd122; b = 8'd95;  #10 
a = 8'd122; b = 8'd96;  #10 
a = 8'd122; b = 8'd97;  #10 
a = 8'd122; b = 8'd98;  #10 
a = 8'd122; b = 8'd99;  #10 
a = 8'd122; b = 8'd100;  #10 
a = 8'd122; b = 8'd101;  #10 
a = 8'd122; b = 8'd102;  #10 
a = 8'd122; b = 8'd103;  #10 
a = 8'd122; b = 8'd104;  #10 
a = 8'd122; b = 8'd105;  #10 
a = 8'd122; b = 8'd106;  #10 
a = 8'd122; b = 8'd107;  #10 
a = 8'd122; b = 8'd108;  #10 
a = 8'd122; b = 8'd109;  #10 
a = 8'd122; b = 8'd110;  #10 
a = 8'd122; b = 8'd111;  #10 
a = 8'd122; b = 8'd112;  #10 
a = 8'd122; b = 8'd113;  #10 
a = 8'd122; b = 8'd114;  #10 
a = 8'd122; b = 8'd115;  #10 
a = 8'd122; b = 8'd116;  #10 
a = 8'd122; b = 8'd117;  #10 
a = 8'd122; b = 8'd118;  #10 
a = 8'd122; b = 8'd119;  #10 
a = 8'd122; b = 8'd120;  #10 
a = 8'd122; b = 8'd121;  #10 
a = 8'd122; b = 8'd122;  #10 
a = 8'd122; b = 8'd123;  #10 
a = 8'd122; b = 8'd124;  #10 
a = 8'd122; b = 8'd125;  #10 
a = 8'd122; b = 8'd126;  #10 
a = 8'd122; b = 8'd127;  #10 
a = 8'd122; b = 8'd128;  #10 
a = 8'd122; b = 8'd129;  #10 
a = 8'd122; b = 8'd130;  #10 
a = 8'd122; b = 8'd131;  #10 
a = 8'd122; b = 8'd132;  #10 
a = 8'd122; b = 8'd133;  #10 
a = 8'd122; b = 8'd134;  #10 
a = 8'd122; b = 8'd135;  #10 
a = 8'd122; b = 8'd136;  #10 
a = 8'd122; b = 8'd137;  #10 
a = 8'd122; b = 8'd138;  #10 
a = 8'd122; b = 8'd139;  #10 
a = 8'd122; b = 8'd140;  #10 
a = 8'd122; b = 8'd141;  #10 
a = 8'd122; b = 8'd142;  #10 
a = 8'd122; b = 8'd143;  #10 
a = 8'd122; b = 8'd144;  #10 
a = 8'd122; b = 8'd145;  #10 
a = 8'd122; b = 8'd146;  #10 
a = 8'd122; b = 8'd147;  #10 
a = 8'd122; b = 8'd148;  #10 
a = 8'd122; b = 8'd149;  #10 
a = 8'd122; b = 8'd150;  #10 
a = 8'd122; b = 8'd151;  #10 
a = 8'd122; b = 8'd152;  #10 
a = 8'd122; b = 8'd153;  #10 
a = 8'd122; b = 8'd154;  #10 
a = 8'd122; b = 8'd155;  #10 
a = 8'd122; b = 8'd156;  #10 
a = 8'd122; b = 8'd157;  #10 
a = 8'd122; b = 8'd158;  #10 
a = 8'd122; b = 8'd159;  #10 
a = 8'd122; b = 8'd160;  #10 
a = 8'd122; b = 8'd161;  #10 
a = 8'd122; b = 8'd162;  #10 
a = 8'd122; b = 8'd163;  #10 
a = 8'd122; b = 8'd164;  #10 
a = 8'd122; b = 8'd165;  #10 
a = 8'd122; b = 8'd166;  #10 
a = 8'd122; b = 8'd167;  #10 
a = 8'd122; b = 8'd168;  #10 
a = 8'd122; b = 8'd169;  #10 
a = 8'd122; b = 8'd170;  #10 
a = 8'd122; b = 8'd171;  #10 
a = 8'd122; b = 8'd172;  #10 
a = 8'd122; b = 8'd173;  #10 
a = 8'd122; b = 8'd174;  #10 
a = 8'd122; b = 8'd175;  #10 
a = 8'd122; b = 8'd176;  #10 
a = 8'd122; b = 8'd177;  #10 
a = 8'd122; b = 8'd178;  #10 
a = 8'd122; b = 8'd179;  #10 
a = 8'd122; b = 8'd180;  #10 
a = 8'd122; b = 8'd181;  #10 
a = 8'd122; b = 8'd182;  #10 
a = 8'd122; b = 8'd183;  #10 
a = 8'd122; b = 8'd184;  #10 
a = 8'd122; b = 8'd185;  #10 
a = 8'd122; b = 8'd186;  #10 
a = 8'd122; b = 8'd187;  #10 
a = 8'd122; b = 8'd188;  #10 
a = 8'd122; b = 8'd189;  #10 
a = 8'd122; b = 8'd190;  #10 
a = 8'd122; b = 8'd191;  #10 
a = 8'd122; b = 8'd192;  #10 
a = 8'd122; b = 8'd193;  #10 
a = 8'd122; b = 8'd194;  #10 
a = 8'd122; b = 8'd195;  #10 
a = 8'd122; b = 8'd196;  #10 
a = 8'd122; b = 8'd197;  #10 
a = 8'd122; b = 8'd198;  #10 
a = 8'd122; b = 8'd199;  #10 
a = 8'd122; b = 8'd200;  #10 
a = 8'd122; b = 8'd201;  #10 
a = 8'd122; b = 8'd202;  #10 
a = 8'd122; b = 8'd203;  #10 
a = 8'd122; b = 8'd204;  #10 
a = 8'd122; b = 8'd205;  #10 
a = 8'd122; b = 8'd206;  #10 
a = 8'd122; b = 8'd207;  #10 
a = 8'd122; b = 8'd208;  #10 
a = 8'd122; b = 8'd209;  #10 
a = 8'd122; b = 8'd210;  #10 
a = 8'd122; b = 8'd211;  #10 
a = 8'd122; b = 8'd212;  #10 
a = 8'd122; b = 8'd213;  #10 
a = 8'd122; b = 8'd214;  #10 
a = 8'd122; b = 8'd215;  #10 
a = 8'd122; b = 8'd216;  #10 
a = 8'd122; b = 8'd217;  #10 
a = 8'd122; b = 8'd218;  #10 
a = 8'd122; b = 8'd219;  #10 
a = 8'd122; b = 8'd220;  #10 
a = 8'd122; b = 8'd221;  #10 
a = 8'd122; b = 8'd222;  #10 
a = 8'd122; b = 8'd223;  #10 
a = 8'd122; b = 8'd224;  #10 
a = 8'd122; b = 8'd225;  #10 
a = 8'd122; b = 8'd226;  #10 
a = 8'd122; b = 8'd227;  #10 
a = 8'd122; b = 8'd228;  #10 
a = 8'd122; b = 8'd229;  #10 
a = 8'd122; b = 8'd230;  #10 
a = 8'd122; b = 8'd231;  #10 
a = 8'd122; b = 8'd232;  #10 
a = 8'd122; b = 8'd233;  #10 
a = 8'd122; b = 8'd234;  #10 
a = 8'd122; b = 8'd235;  #10 
a = 8'd122; b = 8'd236;  #10 
a = 8'd122; b = 8'd237;  #10 
a = 8'd122; b = 8'd238;  #10 
a = 8'd122; b = 8'd239;  #10 
a = 8'd122; b = 8'd240;  #10 
a = 8'd122; b = 8'd241;  #10 
a = 8'd122; b = 8'd242;  #10 
a = 8'd122; b = 8'd243;  #10 
a = 8'd122; b = 8'd244;  #10 
a = 8'd122; b = 8'd245;  #10 
a = 8'd122; b = 8'd246;  #10 
a = 8'd122; b = 8'd247;  #10 
a = 8'd122; b = 8'd248;  #10 
a = 8'd122; b = 8'd249;  #10 
a = 8'd122; b = 8'd250;  #10 
a = 8'd122; b = 8'd251;  #10 
a = 8'd122; b = 8'd252;  #10 
a = 8'd122; b = 8'd253;  #10 
a = 8'd122; b = 8'd254;  #10 
a = 8'd122; b = 8'd255;  #10 
a = 8'd123; b = 8'd0;  #10 
a = 8'd123; b = 8'd1;  #10 
a = 8'd123; b = 8'd2;  #10 
a = 8'd123; b = 8'd3;  #10 
a = 8'd123; b = 8'd4;  #10 
a = 8'd123; b = 8'd5;  #10 
a = 8'd123; b = 8'd6;  #10 
a = 8'd123; b = 8'd7;  #10 
a = 8'd123; b = 8'd8;  #10 
a = 8'd123; b = 8'd9;  #10 
a = 8'd123; b = 8'd10;  #10 
a = 8'd123; b = 8'd11;  #10 
a = 8'd123; b = 8'd12;  #10 
a = 8'd123; b = 8'd13;  #10 
a = 8'd123; b = 8'd14;  #10 
a = 8'd123; b = 8'd15;  #10 
a = 8'd123; b = 8'd16;  #10 
a = 8'd123; b = 8'd17;  #10 
a = 8'd123; b = 8'd18;  #10 
a = 8'd123; b = 8'd19;  #10 
a = 8'd123; b = 8'd20;  #10 
a = 8'd123; b = 8'd21;  #10 
a = 8'd123; b = 8'd22;  #10 
a = 8'd123; b = 8'd23;  #10 
a = 8'd123; b = 8'd24;  #10 
a = 8'd123; b = 8'd25;  #10 
a = 8'd123; b = 8'd26;  #10 
a = 8'd123; b = 8'd27;  #10 
a = 8'd123; b = 8'd28;  #10 
a = 8'd123; b = 8'd29;  #10 
a = 8'd123; b = 8'd30;  #10 
a = 8'd123; b = 8'd31;  #10 
a = 8'd123; b = 8'd32;  #10 
a = 8'd123; b = 8'd33;  #10 
a = 8'd123; b = 8'd34;  #10 
a = 8'd123; b = 8'd35;  #10 
a = 8'd123; b = 8'd36;  #10 
a = 8'd123; b = 8'd37;  #10 
a = 8'd123; b = 8'd38;  #10 
a = 8'd123; b = 8'd39;  #10 
a = 8'd123; b = 8'd40;  #10 
a = 8'd123; b = 8'd41;  #10 
a = 8'd123; b = 8'd42;  #10 
a = 8'd123; b = 8'd43;  #10 
a = 8'd123; b = 8'd44;  #10 
a = 8'd123; b = 8'd45;  #10 
a = 8'd123; b = 8'd46;  #10 
a = 8'd123; b = 8'd47;  #10 
a = 8'd123; b = 8'd48;  #10 
a = 8'd123; b = 8'd49;  #10 
a = 8'd123; b = 8'd50;  #10 
a = 8'd123; b = 8'd51;  #10 
a = 8'd123; b = 8'd52;  #10 
a = 8'd123; b = 8'd53;  #10 
a = 8'd123; b = 8'd54;  #10 
a = 8'd123; b = 8'd55;  #10 
a = 8'd123; b = 8'd56;  #10 
a = 8'd123; b = 8'd57;  #10 
a = 8'd123; b = 8'd58;  #10 
a = 8'd123; b = 8'd59;  #10 
a = 8'd123; b = 8'd60;  #10 
a = 8'd123; b = 8'd61;  #10 
a = 8'd123; b = 8'd62;  #10 
a = 8'd123; b = 8'd63;  #10 
a = 8'd123; b = 8'd64;  #10 
a = 8'd123; b = 8'd65;  #10 
a = 8'd123; b = 8'd66;  #10 
a = 8'd123; b = 8'd67;  #10 
a = 8'd123; b = 8'd68;  #10 
a = 8'd123; b = 8'd69;  #10 
a = 8'd123; b = 8'd70;  #10 
a = 8'd123; b = 8'd71;  #10 
a = 8'd123; b = 8'd72;  #10 
a = 8'd123; b = 8'd73;  #10 
a = 8'd123; b = 8'd74;  #10 
a = 8'd123; b = 8'd75;  #10 
a = 8'd123; b = 8'd76;  #10 
a = 8'd123; b = 8'd77;  #10 
a = 8'd123; b = 8'd78;  #10 
a = 8'd123; b = 8'd79;  #10 
a = 8'd123; b = 8'd80;  #10 
a = 8'd123; b = 8'd81;  #10 
a = 8'd123; b = 8'd82;  #10 
a = 8'd123; b = 8'd83;  #10 
a = 8'd123; b = 8'd84;  #10 
a = 8'd123; b = 8'd85;  #10 
a = 8'd123; b = 8'd86;  #10 
a = 8'd123; b = 8'd87;  #10 
a = 8'd123; b = 8'd88;  #10 
a = 8'd123; b = 8'd89;  #10 
a = 8'd123; b = 8'd90;  #10 
a = 8'd123; b = 8'd91;  #10 
a = 8'd123; b = 8'd92;  #10 
a = 8'd123; b = 8'd93;  #10 
a = 8'd123; b = 8'd94;  #10 
a = 8'd123; b = 8'd95;  #10 
a = 8'd123; b = 8'd96;  #10 
a = 8'd123; b = 8'd97;  #10 
a = 8'd123; b = 8'd98;  #10 
a = 8'd123; b = 8'd99;  #10 
a = 8'd123; b = 8'd100;  #10 
a = 8'd123; b = 8'd101;  #10 
a = 8'd123; b = 8'd102;  #10 
a = 8'd123; b = 8'd103;  #10 
a = 8'd123; b = 8'd104;  #10 
a = 8'd123; b = 8'd105;  #10 
a = 8'd123; b = 8'd106;  #10 
a = 8'd123; b = 8'd107;  #10 
a = 8'd123; b = 8'd108;  #10 
a = 8'd123; b = 8'd109;  #10 
a = 8'd123; b = 8'd110;  #10 
a = 8'd123; b = 8'd111;  #10 
a = 8'd123; b = 8'd112;  #10 
a = 8'd123; b = 8'd113;  #10 
a = 8'd123; b = 8'd114;  #10 
a = 8'd123; b = 8'd115;  #10 
a = 8'd123; b = 8'd116;  #10 
a = 8'd123; b = 8'd117;  #10 
a = 8'd123; b = 8'd118;  #10 
a = 8'd123; b = 8'd119;  #10 
a = 8'd123; b = 8'd120;  #10 
a = 8'd123; b = 8'd121;  #10 
a = 8'd123; b = 8'd122;  #10 
a = 8'd123; b = 8'd123;  #10 
a = 8'd123; b = 8'd124;  #10 
a = 8'd123; b = 8'd125;  #10 
a = 8'd123; b = 8'd126;  #10 
a = 8'd123; b = 8'd127;  #10 
a = 8'd123; b = 8'd128;  #10 
a = 8'd123; b = 8'd129;  #10 
a = 8'd123; b = 8'd130;  #10 
a = 8'd123; b = 8'd131;  #10 
a = 8'd123; b = 8'd132;  #10 
a = 8'd123; b = 8'd133;  #10 
a = 8'd123; b = 8'd134;  #10 
a = 8'd123; b = 8'd135;  #10 
a = 8'd123; b = 8'd136;  #10 
a = 8'd123; b = 8'd137;  #10 
a = 8'd123; b = 8'd138;  #10 
a = 8'd123; b = 8'd139;  #10 
a = 8'd123; b = 8'd140;  #10 
a = 8'd123; b = 8'd141;  #10 
a = 8'd123; b = 8'd142;  #10 
a = 8'd123; b = 8'd143;  #10 
a = 8'd123; b = 8'd144;  #10 
a = 8'd123; b = 8'd145;  #10 
a = 8'd123; b = 8'd146;  #10 
a = 8'd123; b = 8'd147;  #10 
a = 8'd123; b = 8'd148;  #10 
a = 8'd123; b = 8'd149;  #10 
a = 8'd123; b = 8'd150;  #10 
a = 8'd123; b = 8'd151;  #10 
a = 8'd123; b = 8'd152;  #10 
a = 8'd123; b = 8'd153;  #10 
a = 8'd123; b = 8'd154;  #10 
a = 8'd123; b = 8'd155;  #10 
a = 8'd123; b = 8'd156;  #10 
a = 8'd123; b = 8'd157;  #10 
a = 8'd123; b = 8'd158;  #10 
a = 8'd123; b = 8'd159;  #10 
a = 8'd123; b = 8'd160;  #10 
a = 8'd123; b = 8'd161;  #10 
a = 8'd123; b = 8'd162;  #10 
a = 8'd123; b = 8'd163;  #10 
a = 8'd123; b = 8'd164;  #10 
a = 8'd123; b = 8'd165;  #10 
a = 8'd123; b = 8'd166;  #10 
a = 8'd123; b = 8'd167;  #10 
a = 8'd123; b = 8'd168;  #10 
a = 8'd123; b = 8'd169;  #10 
a = 8'd123; b = 8'd170;  #10 
a = 8'd123; b = 8'd171;  #10 
a = 8'd123; b = 8'd172;  #10 
a = 8'd123; b = 8'd173;  #10 
a = 8'd123; b = 8'd174;  #10 
a = 8'd123; b = 8'd175;  #10 
a = 8'd123; b = 8'd176;  #10 
a = 8'd123; b = 8'd177;  #10 
a = 8'd123; b = 8'd178;  #10 
a = 8'd123; b = 8'd179;  #10 
a = 8'd123; b = 8'd180;  #10 
a = 8'd123; b = 8'd181;  #10 
a = 8'd123; b = 8'd182;  #10 
a = 8'd123; b = 8'd183;  #10 
a = 8'd123; b = 8'd184;  #10 
a = 8'd123; b = 8'd185;  #10 
a = 8'd123; b = 8'd186;  #10 
a = 8'd123; b = 8'd187;  #10 
a = 8'd123; b = 8'd188;  #10 
a = 8'd123; b = 8'd189;  #10 
a = 8'd123; b = 8'd190;  #10 
a = 8'd123; b = 8'd191;  #10 
a = 8'd123; b = 8'd192;  #10 
a = 8'd123; b = 8'd193;  #10 
a = 8'd123; b = 8'd194;  #10 
a = 8'd123; b = 8'd195;  #10 
a = 8'd123; b = 8'd196;  #10 
a = 8'd123; b = 8'd197;  #10 
a = 8'd123; b = 8'd198;  #10 
a = 8'd123; b = 8'd199;  #10 
a = 8'd123; b = 8'd200;  #10 
a = 8'd123; b = 8'd201;  #10 
a = 8'd123; b = 8'd202;  #10 
a = 8'd123; b = 8'd203;  #10 
a = 8'd123; b = 8'd204;  #10 
a = 8'd123; b = 8'd205;  #10 
a = 8'd123; b = 8'd206;  #10 
a = 8'd123; b = 8'd207;  #10 
a = 8'd123; b = 8'd208;  #10 
a = 8'd123; b = 8'd209;  #10 
a = 8'd123; b = 8'd210;  #10 
a = 8'd123; b = 8'd211;  #10 
a = 8'd123; b = 8'd212;  #10 
a = 8'd123; b = 8'd213;  #10 
a = 8'd123; b = 8'd214;  #10 
a = 8'd123; b = 8'd215;  #10 
a = 8'd123; b = 8'd216;  #10 
a = 8'd123; b = 8'd217;  #10 
a = 8'd123; b = 8'd218;  #10 
a = 8'd123; b = 8'd219;  #10 
a = 8'd123; b = 8'd220;  #10 
a = 8'd123; b = 8'd221;  #10 
a = 8'd123; b = 8'd222;  #10 
a = 8'd123; b = 8'd223;  #10 
a = 8'd123; b = 8'd224;  #10 
a = 8'd123; b = 8'd225;  #10 
a = 8'd123; b = 8'd226;  #10 
a = 8'd123; b = 8'd227;  #10 
a = 8'd123; b = 8'd228;  #10 
a = 8'd123; b = 8'd229;  #10 
a = 8'd123; b = 8'd230;  #10 
a = 8'd123; b = 8'd231;  #10 
a = 8'd123; b = 8'd232;  #10 
a = 8'd123; b = 8'd233;  #10 
a = 8'd123; b = 8'd234;  #10 
a = 8'd123; b = 8'd235;  #10 
a = 8'd123; b = 8'd236;  #10 
a = 8'd123; b = 8'd237;  #10 
a = 8'd123; b = 8'd238;  #10 
a = 8'd123; b = 8'd239;  #10 
a = 8'd123; b = 8'd240;  #10 
a = 8'd123; b = 8'd241;  #10 
a = 8'd123; b = 8'd242;  #10 
a = 8'd123; b = 8'd243;  #10 
a = 8'd123; b = 8'd244;  #10 
a = 8'd123; b = 8'd245;  #10 
a = 8'd123; b = 8'd246;  #10 
a = 8'd123; b = 8'd247;  #10 
a = 8'd123; b = 8'd248;  #10 
a = 8'd123; b = 8'd249;  #10 
a = 8'd123; b = 8'd250;  #10 
a = 8'd123; b = 8'd251;  #10 
a = 8'd123; b = 8'd252;  #10 
a = 8'd123; b = 8'd253;  #10 
a = 8'd123; b = 8'd254;  #10 
a = 8'd123; b = 8'd255;  #10 
a = 8'd124; b = 8'd0;  #10 
a = 8'd124; b = 8'd1;  #10 
a = 8'd124; b = 8'd2;  #10 
a = 8'd124; b = 8'd3;  #10 
a = 8'd124; b = 8'd4;  #10 
a = 8'd124; b = 8'd5;  #10 
a = 8'd124; b = 8'd6;  #10 
a = 8'd124; b = 8'd7;  #10 
a = 8'd124; b = 8'd8;  #10 
a = 8'd124; b = 8'd9;  #10 
a = 8'd124; b = 8'd10;  #10 
a = 8'd124; b = 8'd11;  #10 
a = 8'd124; b = 8'd12;  #10 
a = 8'd124; b = 8'd13;  #10 
a = 8'd124; b = 8'd14;  #10 
a = 8'd124; b = 8'd15;  #10 
a = 8'd124; b = 8'd16;  #10 
a = 8'd124; b = 8'd17;  #10 
a = 8'd124; b = 8'd18;  #10 
a = 8'd124; b = 8'd19;  #10 
a = 8'd124; b = 8'd20;  #10 
a = 8'd124; b = 8'd21;  #10 
a = 8'd124; b = 8'd22;  #10 
a = 8'd124; b = 8'd23;  #10 
a = 8'd124; b = 8'd24;  #10 
a = 8'd124; b = 8'd25;  #10 
a = 8'd124; b = 8'd26;  #10 
a = 8'd124; b = 8'd27;  #10 
a = 8'd124; b = 8'd28;  #10 
a = 8'd124; b = 8'd29;  #10 
a = 8'd124; b = 8'd30;  #10 
a = 8'd124; b = 8'd31;  #10 
a = 8'd124; b = 8'd32;  #10 
a = 8'd124; b = 8'd33;  #10 
a = 8'd124; b = 8'd34;  #10 
a = 8'd124; b = 8'd35;  #10 
a = 8'd124; b = 8'd36;  #10 
a = 8'd124; b = 8'd37;  #10 
a = 8'd124; b = 8'd38;  #10 
a = 8'd124; b = 8'd39;  #10 
a = 8'd124; b = 8'd40;  #10 
a = 8'd124; b = 8'd41;  #10 
a = 8'd124; b = 8'd42;  #10 
a = 8'd124; b = 8'd43;  #10 
a = 8'd124; b = 8'd44;  #10 
a = 8'd124; b = 8'd45;  #10 
a = 8'd124; b = 8'd46;  #10 
a = 8'd124; b = 8'd47;  #10 
a = 8'd124; b = 8'd48;  #10 
a = 8'd124; b = 8'd49;  #10 
a = 8'd124; b = 8'd50;  #10 
a = 8'd124; b = 8'd51;  #10 
a = 8'd124; b = 8'd52;  #10 
a = 8'd124; b = 8'd53;  #10 
a = 8'd124; b = 8'd54;  #10 
a = 8'd124; b = 8'd55;  #10 
a = 8'd124; b = 8'd56;  #10 
a = 8'd124; b = 8'd57;  #10 
a = 8'd124; b = 8'd58;  #10 
a = 8'd124; b = 8'd59;  #10 
a = 8'd124; b = 8'd60;  #10 
a = 8'd124; b = 8'd61;  #10 
a = 8'd124; b = 8'd62;  #10 
a = 8'd124; b = 8'd63;  #10 
a = 8'd124; b = 8'd64;  #10 
a = 8'd124; b = 8'd65;  #10 
a = 8'd124; b = 8'd66;  #10 
a = 8'd124; b = 8'd67;  #10 
a = 8'd124; b = 8'd68;  #10 
a = 8'd124; b = 8'd69;  #10 
a = 8'd124; b = 8'd70;  #10 
a = 8'd124; b = 8'd71;  #10 
a = 8'd124; b = 8'd72;  #10 
a = 8'd124; b = 8'd73;  #10 
a = 8'd124; b = 8'd74;  #10 
a = 8'd124; b = 8'd75;  #10 
a = 8'd124; b = 8'd76;  #10 
a = 8'd124; b = 8'd77;  #10 
a = 8'd124; b = 8'd78;  #10 
a = 8'd124; b = 8'd79;  #10 
a = 8'd124; b = 8'd80;  #10 
a = 8'd124; b = 8'd81;  #10 
a = 8'd124; b = 8'd82;  #10 
a = 8'd124; b = 8'd83;  #10 
a = 8'd124; b = 8'd84;  #10 
a = 8'd124; b = 8'd85;  #10 
a = 8'd124; b = 8'd86;  #10 
a = 8'd124; b = 8'd87;  #10 
a = 8'd124; b = 8'd88;  #10 
a = 8'd124; b = 8'd89;  #10 
a = 8'd124; b = 8'd90;  #10 
a = 8'd124; b = 8'd91;  #10 
a = 8'd124; b = 8'd92;  #10 
a = 8'd124; b = 8'd93;  #10 
a = 8'd124; b = 8'd94;  #10 
a = 8'd124; b = 8'd95;  #10 
a = 8'd124; b = 8'd96;  #10 
a = 8'd124; b = 8'd97;  #10 
a = 8'd124; b = 8'd98;  #10 
a = 8'd124; b = 8'd99;  #10 
a = 8'd124; b = 8'd100;  #10 
a = 8'd124; b = 8'd101;  #10 
a = 8'd124; b = 8'd102;  #10 
a = 8'd124; b = 8'd103;  #10 
a = 8'd124; b = 8'd104;  #10 
a = 8'd124; b = 8'd105;  #10 
a = 8'd124; b = 8'd106;  #10 
a = 8'd124; b = 8'd107;  #10 
a = 8'd124; b = 8'd108;  #10 
a = 8'd124; b = 8'd109;  #10 
a = 8'd124; b = 8'd110;  #10 
a = 8'd124; b = 8'd111;  #10 
a = 8'd124; b = 8'd112;  #10 
a = 8'd124; b = 8'd113;  #10 
a = 8'd124; b = 8'd114;  #10 
a = 8'd124; b = 8'd115;  #10 
a = 8'd124; b = 8'd116;  #10 
a = 8'd124; b = 8'd117;  #10 
a = 8'd124; b = 8'd118;  #10 
a = 8'd124; b = 8'd119;  #10 
a = 8'd124; b = 8'd120;  #10 
a = 8'd124; b = 8'd121;  #10 
a = 8'd124; b = 8'd122;  #10 
a = 8'd124; b = 8'd123;  #10 
a = 8'd124; b = 8'd124;  #10 
a = 8'd124; b = 8'd125;  #10 
a = 8'd124; b = 8'd126;  #10 
a = 8'd124; b = 8'd127;  #10 
a = 8'd124; b = 8'd128;  #10 
a = 8'd124; b = 8'd129;  #10 
a = 8'd124; b = 8'd130;  #10 
a = 8'd124; b = 8'd131;  #10 
a = 8'd124; b = 8'd132;  #10 
a = 8'd124; b = 8'd133;  #10 
a = 8'd124; b = 8'd134;  #10 
a = 8'd124; b = 8'd135;  #10 
a = 8'd124; b = 8'd136;  #10 
a = 8'd124; b = 8'd137;  #10 
a = 8'd124; b = 8'd138;  #10 
a = 8'd124; b = 8'd139;  #10 
a = 8'd124; b = 8'd140;  #10 
a = 8'd124; b = 8'd141;  #10 
a = 8'd124; b = 8'd142;  #10 
a = 8'd124; b = 8'd143;  #10 
a = 8'd124; b = 8'd144;  #10 
a = 8'd124; b = 8'd145;  #10 
a = 8'd124; b = 8'd146;  #10 
a = 8'd124; b = 8'd147;  #10 
a = 8'd124; b = 8'd148;  #10 
a = 8'd124; b = 8'd149;  #10 
a = 8'd124; b = 8'd150;  #10 
a = 8'd124; b = 8'd151;  #10 
a = 8'd124; b = 8'd152;  #10 
a = 8'd124; b = 8'd153;  #10 
a = 8'd124; b = 8'd154;  #10 
a = 8'd124; b = 8'd155;  #10 
a = 8'd124; b = 8'd156;  #10 
a = 8'd124; b = 8'd157;  #10 
a = 8'd124; b = 8'd158;  #10 
a = 8'd124; b = 8'd159;  #10 
a = 8'd124; b = 8'd160;  #10 
a = 8'd124; b = 8'd161;  #10 
a = 8'd124; b = 8'd162;  #10 
a = 8'd124; b = 8'd163;  #10 
a = 8'd124; b = 8'd164;  #10 
a = 8'd124; b = 8'd165;  #10 
a = 8'd124; b = 8'd166;  #10 
a = 8'd124; b = 8'd167;  #10 
a = 8'd124; b = 8'd168;  #10 
a = 8'd124; b = 8'd169;  #10 
a = 8'd124; b = 8'd170;  #10 
a = 8'd124; b = 8'd171;  #10 
a = 8'd124; b = 8'd172;  #10 
a = 8'd124; b = 8'd173;  #10 
a = 8'd124; b = 8'd174;  #10 
a = 8'd124; b = 8'd175;  #10 
a = 8'd124; b = 8'd176;  #10 
a = 8'd124; b = 8'd177;  #10 
a = 8'd124; b = 8'd178;  #10 
a = 8'd124; b = 8'd179;  #10 
a = 8'd124; b = 8'd180;  #10 
a = 8'd124; b = 8'd181;  #10 
a = 8'd124; b = 8'd182;  #10 
a = 8'd124; b = 8'd183;  #10 
a = 8'd124; b = 8'd184;  #10 
a = 8'd124; b = 8'd185;  #10 
a = 8'd124; b = 8'd186;  #10 
a = 8'd124; b = 8'd187;  #10 
a = 8'd124; b = 8'd188;  #10 
a = 8'd124; b = 8'd189;  #10 
a = 8'd124; b = 8'd190;  #10 
a = 8'd124; b = 8'd191;  #10 
a = 8'd124; b = 8'd192;  #10 
a = 8'd124; b = 8'd193;  #10 
a = 8'd124; b = 8'd194;  #10 
a = 8'd124; b = 8'd195;  #10 
a = 8'd124; b = 8'd196;  #10 
a = 8'd124; b = 8'd197;  #10 
a = 8'd124; b = 8'd198;  #10 
a = 8'd124; b = 8'd199;  #10 
a = 8'd124; b = 8'd200;  #10 
a = 8'd124; b = 8'd201;  #10 
a = 8'd124; b = 8'd202;  #10 
a = 8'd124; b = 8'd203;  #10 
a = 8'd124; b = 8'd204;  #10 
a = 8'd124; b = 8'd205;  #10 
a = 8'd124; b = 8'd206;  #10 
a = 8'd124; b = 8'd207;  #10 
a = 8'd124; b = 8'd208;  #10 
a = 8'd124; b = 8'd209;  #10 
a = 8'd124; b = 8'd210;  #10 
a = 8'd124; b = 8'd211;  #10 
a = 8'd124; b = 8'd212;  #10 
a = 8'd124; b = 8'd213;  #10 
a = 8'd124; b = 8'd214;  #10 
a = 8'd124; b = 8'd215;  #10 
a = 8'd124; b = 8'd216;  #10 
a = 8'd124; b = 8'd217;  #10 
a = 8'd124; b = 8'd218;  #10 
a = 8'd124; b = 8'd219;  #10 
a = 8'd124; b = 8'd220;  #10 
a = 8'd124; b = 8'd221;  #10 
a = 8'd124; b = 8'd222;  #10 
a = 8'd124; b = 8'd223;  #10 
a = 8'd124; b = 8'd224;  #10 
a = 8'd124; b = 8'd225;  #10 
a = 8'd124; b = 8'd226;  #10 
a = 8'd124; b = 8'd227;  #10 
a = 8'd124; b = 8'd228;  #10 
a = 8'd124; b = 8'd229;  #10 
a = 8'd124; b = 8'd230;  #10 
a = 8'd124; b = 8'd231;  #10 
a = 8'd124; b = 8'd232;  #10 
a = 8'd124; b = 8'd233;  #10 
a = 8'd124; b = 8'd234;  #10 
a = 8'd124; b = 8'd235;  #10 
a = 8'd124; b = 8'd236;  #10 
a = 8'd124; b = 8'd237;  #10 
a = 8'd124; b = 8'd238;  #10 
a = 8'd124; b = 8'd239;  #10 
a = 8'd124; b = 8'd240;  #10 
a = 8'd124; b = 8'd241;  #10 
a = 8'd124; b = 8'd242;  #10 
a = 8'd124; b = 8'd243;  #10 
a = 8'd124; b = 8'd244;  #10 
a = 8'd124; b = 8'd245;  #10 
a = 8'd124; b = 8'd246;  #10 
a = 8'd124; b = 8'd247;  #10 
a = 8'd124; b = 8'd248;  #10 
a = 8'd124; b = 8'd249;  #10 
a = 8'd124; b = 8'd250;  #10 
a = 8'd124; b = 8'd251;  #10 
a = 8'd124; b = 8'd252;  #10 
a = 8'd124; b = 8'd253;  #10 
a = 8'd124; b = 8'd254;  #10 
a = 8'd124; b = 8'd255;  #10 
a = 8'd125; b = 8'd0;  #10 
a = 8'd125; b = 8'd1;  #10 
a = 8'd125; b = 8'd2;  #10 
a = 8'd125; b = 8'd3;  #10 
a = 8'd125; b = 8'd4;  #10 
a = 8'd125; b = 8'd5;  #10 
a = 8'd125; b = 8'd6;  #10 
a = 8'd125; b = 8'd7;  #10 
a = 8'd125; b = 8'd8;  #10 
a = 8'd125; b = 8'd9;  #10 
a = 8'd125; b = 8'd10;  #10 
a = 8'd125; b = 8'd11;  #10 
a = 8'd125; b = 8'd12;  #10 
a = 8'd125; b = 8'd13;  #10 
a = 8'd125; b = 8'd14;  #10 
a = 8'd125; b = 8'd15;  #10 
a = 8'd125; b = 8'd16;  #10 
a = 8'd125; b = 8'd17;  #10 
a = 8'd125; b = 8'd18;  #10 
a = 8'd125; b = 8'd19;  #10 
a = 8'd125; b = 8'd20;  #10 
a = 8'd125; b = 8'd21;  #10 
a = 8'd125; b = 8'd22;  #10 
a = 8'd125; b = 8'd23;  #10 
a = 8'd125; b = 8'd24;  #10 
a = 8'd125; b = 8'd25;  #10 
a = 8'd125; b = 8'd26;  #10 
a = 8'd125; b = 8'd27;  #10 
a = 8'd125; b = 8'd28;  #10 
a = 8'd125; b = 8'd29;  #10 
a = 8'd125; b = 8'd30;  #10 
a = 8'd125; b = 8'd31;  #10 
a = 8'd125; b = 8'd32;  #10 
a = 8'd125; b = 8'd33;  #10 
a = 8'd125; b = 8'd34;  #10 
a = 8'd125; b = 8'd35;  #10 
a = 8'd125; b = 8'd36;  #10 
a = 8'd125; b = 8'd37;  #10 
a = 8'd125; b = 8'd38;  #10 
a = 8'd125; b = 8'd39;  #10 
a = 8'd125; b = 8'd40;  #10 
a = 8'd125; b = 8'd41;  #10 
a = 8'd125; b = 8'd42;  #10 
a = 8'd125; b = 8'd43;  #10 
a = 8'd125; b = 8'd44;  #10 
a = 8'd125; b = 8'd45;  #10 
a = 8'd125; b = 8'd46;  #10 
a = 8'd125; b = 8'd47;  #10 
a = 8'd125; b = 8'd48;  #10 
a = 8'd125; b = 8'd49;  #10 
a = 8'd125; b = 8'd50;  #10 
a = 8'd125; b = 8'd51;  #10 
a = 8'd125; b = 8'd52;  #10 
a = 8'd125; b = 8'd53;  #10 
a = 8'd125; b = 8'd54;  #10 
a = 8'd125; b = 8'd55;  #10 
a = 8'd125; b = 8'd56;  #10 
a = 8'd125; b = 8'd57;  #10 
a = 8'd125; b = 8'd58;  #10 
a = 8'd125; b = 8'd59;  #10 
a = 8'd125; b = 8'd60;  #10 
a = 8'd125; b = 8'd61;  #10 
a = 8'd125; b = 8'd62;  #10 
a = 8'd125; b = 8'd63;  #10 
a = 8'd125; b = 8'd64;  #10 
a = 8'd125; b = 8'd65;  #10 
a = 8'd125; b = 8'd66;  #10 
a = 8'd125; b = 8'd67;  #10 
a = 8'd125; b = 8'd68;  #10 
a = 8'd125; b = 8'd69;  #10 
a = 8'd125; b = 8'd70;  #10 
a = 8'd125; b = 8'd71;  #10 
a = 8'd125; b = 8'd72;  #10 
a = 8'd125; b = 8'd73;  #10 
a = 8'd125; b = 8'd74;  #10 
a = 8'd125; b = 8'd75;  #10 
a = 8'd125; b = 8'd76;  #10 
a = 8'd125; b = 8'd77;  #10 
a = 8'd125; b = 8'd78;  #10 
a = 8'd125; b = 8'd79;  #10 
a = 8'd125; b = 8'd80;  #10 
a = 8'd125; b = 8'd81;  #10 
a = 8'd125; b = 8'd82;  #10 
a = 8'd125; b = 8'd83;  #10 
a = 8'd125; b = 8'd84;  #10 
a = 8'd125; b = 8'd85;  #10 
a = 8'd125; b = 8'd86;  #10 
a = 8'd125; b = 8'd87;  #10 
a = 8'd125; b = 8'd88;  #10 
a = 8'd125; b = 8'd89;  #10 
a = 8'd125; b = 8'd90;  #10 
a = 8'd125; b = 8'd91;  #10 
a = 8'd125; b = 8'd92;  #10 
a = 8'd125; b = 8'd93;  #10 
a = 8'd125; b = 8'd94;  #10 
a = 8'd125; b = 8'd95;  #10 
a = 8'd125; b = 8'd96;  #10 
a = 8'd125; b = 8'd97;  #10 
a = 8'd125; b = 8'd98;  #10 
a = 8'd125; b = 8'd99;  #10 
a = 8'd125; b = 8'd100;  #10 
a = 8'd125; b = 8'd101;  #10 
a = 8'd125; b = 8'd102;  #10 
a = 8'd125; b = 8'd103;  #10 
a = 8'd125; b = 8'd104;  #10 
a = 8'd125; b = 8'd105;  #10 
a = 8'd125; b = 8'd106;  #10 
a = 8'd125; b = 8'd107;  #10 
a = 8'd125; b = 8'd108;  #10 
a = 8'd125; b = 8'd109;  #10 
a = 8'd125; b = 8'd110;  #10 
a = 8'd125; b = 8'd111;  #10 
a = 8'd125; b = 8'd112;  #10 
a = 8'd125; b = 8'd113;  #10 
a = 8'd125; b = 8'd114;  #10 
a = 8'd125; b = 8'd115;  #10 
a = 8'd125; b = 8'd116;  #10 
a = 8'd125; b = 8'd117;  #10 
a = 8'd125; b = 8'd118;  #10 
a = 8'd125; b = 8'd119;  #10 
a = 8'd125; b = 8'd120;  #10 
a = 8'd125; b = 8'd121;  #10 
a = 8'd125; b = 8'd122;  #10 
a = 8'd125; b = 8'd123;  #10 
a = 8'd125; b = 8'd124;  #10 
a = 8'd125; b = 8'd125;  #10 
a = 8'd125; b = 8'd126;  #10 
a = 8'd125; b = 8'd127;  #10 
a = 8'd125; b = 8'd128;  #10 
a = 8'd125; b = 8'd129;  #10 
a = 8'd125; b = 8'd130;  #10 
a = 8'd125; b = 8'd131;  #10 
a = 8'd125; b = 8'd132;  #10 
a = 8'd125; b = 8'd133;  #10 
a = 8'd125; b = 8'd134;  #10 
a = 8'd125; b = 8'd135;  #10 
a = 8'd125; b = 8'd136;  #10 
a = 8'd125; b = 8'd137;  #10 
a = 8'd125; b = 8'd138;  #10 
a = 8'd125; b = 8'd139;  #10 
a = 8'd125; b = 8'd140;  #10 
a = 8'd125; b = 8'd141;  #10 
a = 8'd125; b = 8'd142;  #10 
a = 8'd125; b = 8'd143;  #10 
a = 8'd125; b = 8'd144;  #10 
a = 8'd125; b = 8'd145;  #10 
a = 8'd125; b = 8'd146;  #10 
a = 8'd125; b = 8'd147;  #10 
a = 8'd125; b = 8'd148;  #10 
a = 8'd125; b = 8'd149;  #10 
a = 8'd125; b = 8'd150;  #10 
a = 8'd125; b = 8'd151;  #10 
a = 8'd125; b = 8'd152;  #10 
a = 8'd125; b = 8'd153;  #10 
a = 8'd125; b = 8'd154;  #10 
a = 8'd125; b = 8'd155;  #10 
a = 8'd125; b = 8'd156;  #10 
a = 8'd125; b = 8'd157;  #10 
a = 8'd125; b = 8'd158;  #10 
a = 8'd125; b = 8'd159;  #10 
a = 8'd125; b = 8'd160;  #10 
a = 8'd125; b = 8'd161;  #10 
a = 8'd125; b = 8'd162;  #10 
a = 8'd125; b = 8'd163;  #10 
a = 8'd125; b = 8'd164;  #10 
a = 8'd125; b = 8'd165;  #10 
a = 8'd125; b = 8'd166;  #10 
a = 8'd125; b = 8'd167;  #10 
a = 8'd125; b = 8'd168;  #10 
a = 8'd125; b = 8'd169;  #10 
a = 8'd125; b = 8'd170;  #10 
a = 8'd125; b = 8'd171;  #10 
a = 8'd125; b = 8'd172;  #10 
a = 8'd125; b = 8'd173;  #10 
a = 8'd125; b = 8'd174;  #10 
a = 8'd125; b = 8'd175;  #10 
a = 8'd125; b = 8'd176;  #10 
a = 8'd125; b = 8'd177;  #10 
a = 8'd125; b = 8'd178;  #10 
a = 8'd125; b = 8'd179;  #10 
a = 8'd125; b = 8'd180;  #10 
a = 8'd125; b = 8'd181;  #10 
a = 8'd125; b = 8'd182;  #10 
a = 8'd125; b = 8'd183;  #10 
a = 8'd125; b = 8'd184;  #10 
a = 8'd125; b = 8'd185;  #10 
a = 8'd125; b = 8'd186;  #10 
a = 8'd125; b = 8'd187;  #10 
a = 8'd125; b = 8'd188;  #10 
a = 8'd125; b = 8'd189;  #10 
a = 8'd125; b = 8'd190;  #10 
a = 8'd125; b = 8'd191;  #10 
a = 8'd125; b = 8'd192;  #10 
a = 8'd125; b = 8'd193;  #10 
a = 8'd125; b = 8'd194;  #10 
a = 8'd125; b = 8'd195;  #10 
a = 8'd125; b = 8'd196;  #10 
a = 8'd125; b = 8'd197;  #10 
a = 8'd125; b = 8'd198;  #10 
a = 8'd125; b = 8'd199;  #10 
a = 8'd125; b = 8'd200;  #10 
a = 8'd125; b = 8'd201;  #10 
a = 8'd125; b = 8'd202;  #10 
a = 8'd125; b = 8'd203;  #10 
a = 8'd125; b = 8'd204;  #10 
a = 8'd125; b = 8'd205;  #10 
a = 8'd125; b = 8'd206;  #10 
a = 8'd125; b = 8'd207;  #10 
a = 8'd125; b = 8'd208;  #10 
a = 8'd125; b = 8'd209;  #10 
a = 8'd125; b = 8'd210;  #10 
a = 8'd125; b = 8'd211;  #10 
a = 8'd125; b = 8'd212;  #10 
a = 8'd125; b = 8'd213;  #10 
a = 8'd125; b = 8'd214;  #10 
a = 8'd125; b = 8'd215;  #10 
a = 8'd125; b = 8'd216;  #10 
a = 8'd125; b = 8'd217;  #10 
a = 8'd125; b = 8'd218;  #10 
a = 8'd125; b = 8'd219;  #10 
a = 8'd125; b = 8'd220;  #10 
a = 8'd125; b = 8'd221;  #10 
a = 8'd125; b = 8'd222;  #10 
a = 8'd125; b = 8'd223;  #10 
a = 8'd125; b = 8'd224;  #10 
a = 8'd125; b = 8'd225;  #10 
a = 8'd125; b = 8'd226;  #10 
a = 8'd125; b = 8'd227;  #10 
a = 8'd125; b = 8'd228;  #10 
a = 8'd125; b = 8'd229;  #10 
a = 8'd125; b = 8'd230;  #10 
a = 8'd125; b = 8'd231;  #10 
a = 8'd125; b = 8'd232;  #10 
a = 8'd125; b = 8'd233;  #10 
a = 8'd125; b = 8'd234;  #10 
a = 8'd125; b = 8'd235;  #10 
a = 8'd125; b = 8'd236;  #10 
a = 8'd125; b = 8'd237;  #10 
a = 8'd125; b = 8'd238;  #10 
a = 8'd125; b = 8'd239;  #10 
a = 8'd125; b = 8'd240;  #10 
a = 8'd125; b = 8'd241;  #10 
a = 8'd125; b = 8'd242;  #10 
a = 8'd125; b = 8'd243;  #10 
a = 8'd125; b = 8'd244;  #10 
a = 8'd125; b = 8'd245;  #10 
a = 8'd125; b = 8'd246;  #10 
a = 8'd125; b = 8'd247;  #10 
a = 8'd125; b = 8'd248;  #10 
a = 8'd125; b = 8'd249;  #10 
a = 8'd125; b = 8'd250;  #10 
a = 8'd125; b = 8'd251;  #10 
a = 8'd125; b = 8'd252;  #10 
a = 8'd125; b = 8'd253;  #10 
a = 8'd125; b = 8'd254;  #10 
a = 8'd125; b = 8'd255;  #10 
a = 8'd126; b = 8'd0;  #10 
a = 8'd126; b = 8'd1;  #10 
a = 8'd126; b = 8'd2;  #10 
a = 8'd126; b = 8'd3;  #10 
a = 8'd126; b = 8'd4;  #10 
a = 8'd126; b = 8'd5;  #10 
a = 8'd126; b = 8'd6;  #10 
a = 8'd126; b = 8'd7;  #10 
a = 8'd126; b = 8'd8;  #10 
a = 8'd126; b = 8'd9;  #10 
a = 8'd126; b = 8'd10;  #10 
a = 8'd126; b = 8'd11;  #10 
a = 8'd126; b = 8'd12;  #10 
a = 8'd126; b = 8'd13;  #10 
a = 8'd126; b = 8'd14;  #10 
a = 8'd126; b = 8'd15;  #10 
a = 8'd126; b = 8'd16;  #10 
a = 8'd126; b = 8'd17;  #10 
a = 8'd126; b = 8'd18;  #10 
a = 8'd126; b = 8'd19;  #10 
a = 8'd126; b = 8'd20;  #10 
a = 8'd126; b = 8'd21;  #10 
a = 8'd126; b = 8'd22;  #10 
a = 8'd126; b = 8'd23;  #10 
a = 8'd126; b = 8'd24;  #10 
a = 8'd126; b = 8'd25;  #10 
a = 8'd126; b = 8'd26;  #10 
a = 8'd126; b = 8'd27;  #10 
a = 8'd126; b = 8'd28;  #10 
a = 8'd126; b = 8'd29;  #10 
a = 8'd126; b = 8'd30;  #10 
a = 8'd126; b = 8'd31;  #10 
a = 8'd126; b = 8'd32;  #10 
a = 8'd126; b = 8'd33;  #10 
a = 8'd126; b = 8'd34;  #10 
a = 8'd126; b = 8'd35;  #10 
a = 8'd126; b = 8'd36;  #10 
a = 8'd126; b = 8'd37;  #10 
a = 8'd126; b = 8'd38;  #10 
a = 8'd126; b = 8'd39;  #10 
a = 8'd126; b = 8'd40;  #10 
a = 8'd126; b = 8'd41;  #10 
a = 8'd126; b = 8'd42;  #10 
a = 8'd126; b = 8'd43;  #10 
a = 8'd126; b = 8'd44;  #10 
a = 8'd126; b = 8'd45;  #10 
a = 8'd126; b = 8'd46;  #10 
a = 8'd126; b = 8'd47;  #10 
a = 8'd126; b = 8'd48;  #10 
a = 8'd126; b = 8'd49;  #10 
a = 8'd126; b = 8'd50;  #10 
a = 8'd126; b = 8'd51;  #10 
a = 8'd126; b = 8'd52;  #10 
a = 8'd126; b = 8'd53;  #10 
a = 8'd126; b = 8'd54;  #10 
a = 8'd126; b = 8'd55;  #10 
a = 8'd126; b = 8'd56;  #10 
a = 8'd126; b = 8'd57;  #10 
a = 8'd126; b = 8'd58;  #10 
a = 8'd126; b = 8'd59;  #10 
a = 8'd126; b = 8'd60;  #10 
a = 8'd126; b = 8'd61;  #10 
a = 8'd126; b = 8'd62;  #10 
a = 8'd126; b = 8'd63;  #10 
a = 8'd126; b = 8'd64;  #10 
a = 8'd126; b = 8'd65;  #10 
a = 8'd126; b = 8'd66;  #10 
a = 8'd126; b = 8'd67;  #10 
a = 8'd126; b = 8'd68;  #10 
a = 8'd126; b = 8'd69;  #10 
a = 8'd126; b = 8'd70;  #10 
a = 8'd126; b = 8'd71;  #10 
a = 8'd126; b = 8'd72;  #10 
a = 8'd126; b = 8'd73;  #10 
a = 8'd126; b = 8'd74;  #10 
a = 8'd126; b = 8'd75;  #10 
a = 8'd126; b = 8'd76;  #10 
a = 8'd126; b = 8'd77;  #10 
a = 8'd126; b = 8'd78;  #10 
a = 8'd126; b = 8'd79;  #10 
a = 8'd126; b = 8'd80;  #10 
a = 8'd126; b = 8'd81;  #10 
a = 8'd126; b = 8'd82;  #10 
a = 8'd126; b = 8'd83;  #10 
a = 8'd126; b = 8'd84;  #10 
a = 8'd126; b = 8'd85;  #10 
a = 8'd126; b = 8'd86;  #10 
a = 8'd126; b = 8'd87;  #10 
a = 8'd126; b = 8'd88;  #10 
a = 8'd126; b = 8'd89;  #10 
a = 8'd126; b = 8'd90;  #10 
a = 8'd126; b = 8'd91;  #10 
a = 8'd126; b = 8'd92;  #10 
a = 8'd126; b = 8'd93;  #10 
a = 8'd126; b = 8'd94;  #10 
a = 8'd126; b = 8'd95;  #10 
a = 8'd126; b = 8'd96;  #10 
a = 8'd126; b = 8'd97;  #10 
a = 8'd126; b = 8'd98;  #10 
a = 8'd126; b = 8'd99;  #10 
a = 8'd126; b = 8'd100;  #10 
a = 8'd126; b = 8'd101;  #10 
a = 8'd126; b = 8'd102;  #10 
a = 8'd126; b = 8'd103;  #10 
a = 8'd126; b = 8'd104;  #10 
a = 8'd126; b = 8'd105;  #10 
a = 8'd126; b = 8'd106;  #10 
a = 8'd126; b = 8'd107;  #10 
a = 8'd126; b = 8'd108;  #10 
a = 8'd126; b = 8'd109;  #10 
a = 8'd126; b = 8'd110;  #10 
a = 8'd126; b = 8'd111;  #10 
a = 8'd126; b = 8'd112;  #10 
a = 8'd126; b = 8'd113;  #10 
a = 8'd126; b = 8'd114;  #10 
a = 8'd126; b = 8'd115;  #10 
a = 8'd126; b = 8'd116;  #10 
a = 8'd126; b = 8'd117;  #10 
a = 8'd126; b = 8'd118;  #10 
a = 8'd126; b = 8'd119;  #10 
a = 8'd126; b = 8'd120;  #10 
a = 8'd126; b = 8'd121;  #10 
a = 8'd126; b = 8'd122;  #10 
a = 8'd126; b = 8'd123;  #10 
a = 8'd126; b = 8'd124;  #10 
a = 8'd126; b = 8'd125;  #10 
a = 8'd126; b = 8'd126;  #10 
a = 8'd126; b = 8'd127;  #10 
a = 8'd126; b = 8'd128;  #10 
a = 8'd126; b = 8'd129;  #10 
a = 8'd126; b = 8'd130;  #10 
a = 8'd126; b = 8'd131;  #10 
a = 8'd126; b = 8'd132;  #10 
a = 8'd126; b = 8'd133;  #10 
a = 8'd126; b = 8'd134;  #10 
a = 8'd126; b = 8'd135;  #10 
a = 8'd126; b = 8'd136;  #10 
a = 8'd126; b = 8'd137;  #10 
a = 8'd126; b = 8'd138;  #10 
a = 8'd126; b = 8'd139;  #10 
a = 8'd126; b = 8'd140;  #10 
a = 8'd126; b = 8'd141;  #10 
a = 8'd126; b = 8'd142;  #10 
a = 8'd126; b = 8'd143;  #10 
a = 8'd126; b = 8'd144;  #10 
a = 8'd126; b = 8'd145;  #10 
a = 8'd126; b = 8'd146;  #10 
a = 8'd126; b = 8'd147;  #10 
a = 8'd126; b = 8'd148;  #10 
a = 8'd126; b = 8'd149;  #10 
a = 8'd126; b = 8'd150;  #10 
a = 8'd126; b = 8'd151;  #10 
a = 8'd126; b = 8'd152;  #10 
a = 8'd126; b = 8'd153;  #10 
a = 8'd126; b = 8'd154;  #10 
a = 8'd126; b = 8'd155;  #10 
a = 8'd126; b = 8'd156;  #10 
a = 8'd126; b = 8'd157;  #10 
a = 8'd126; b = 8'd158;  #10 
a = 8'd126; b = 8'd159;  #10 
a = 8'd126; b = 8'd160;  #10 
a = 8'd126; b = 8'd161;  #10 
a = 8'd126; b = 8'd162;  #10 
a = 8'd126; b = 8'd163;  #10 
a = 8'd126; b = 8'd164;  #10 
a = 8'd126; b = 8'd165;  #10 
a = 8'd126; b = 8'd166;  #10 
a = 8'd126; b = 8'd167;  #10 
a = 8'd126; b = 8'd168;  #10 
a = 8'd126; b = 8'd169;  #10 
a = 8'd126; b = 8'd170;  #10 
a = 8'd126; b = 8'd171;  #10 
a = 8'd126; b = 8'd172;  #10 
a = 8'd126; b = 8'd173;  #10 
a = 8'd126; b = 8'd174;  #10 
a = 8'd126; b = 8'd175;  #10 
a = 8'd126; b = 8'd176;  #10 
a = 8'd126; b = 8'd177;  #10 
a = 8'd126; b = 8'd178;  #10 
a = 8'd126; b = 8'd179;  #10 
a = 8'd126; b = 8'd180;  #10 
a = 8'd126; b = 8'd181;  #10 
a = 8'd126; b = 8'd182;  #10 
a = 8'd126; b = 8'd183;  #10 
a = 8'd126; b = 8'd184;  #10 
a = 8'd126; b = 8'd185;  #10 
a = 8'd126; b = 8'd186;  #10 
a = 8'd126; b = 8'd187;  #10 
a = 8'd126; b = 8'd188;  #10 
a = 8'd126; b = 8'd189;  #10 
a = 8'd126; b = 8'd190;  #10 
a = 8'd126; b = 8'd191;  #10 
a = 8'd126; b = 8'd192;  #10 
a = 8'd126; b = 8'd193;  #10 
a = 8'd126; b = 8'd194;  #10 
a = 8'd126; b = 8'd195;  #10 
a = 8'd126; b = 8'd196;  #10 
a = 8'd126; b = 8'd197;  #10 
a = 8'd126; b = 8'd198;  #10 
a = 8'd126; b = 8'd199;  #10 
a = 8'd126; b = 8'd200;  #10 
a = 8'd126; b = 8'd201;  #10 
a = 8'd126; b = 8'd202;  #10 
a = 8'd126; b = 8'd203;  #10 
a = 8'd126; b = 8'd204;  #10 
a = 8'd126; b = 8'd205;  #10 
a = 8'd126; b = 8'd206;  #10 
a = 8'd126; b = 8'd207;  #10 
a = 8'd126; b = 8'd208;  #10 
a = 8'd126; b = 8'd209;  #10 
a = 8'd126; b = 8'd210;  #10 
a = 8'd126; b = 8'd211;  #10 
a = 8'd126; b = 8'd212;  #10 
a = 8'd126; b = 8'd213;  #10 
a = 8'd126; b = 8'd214;  #10 
a = 8'd126; b = 8'd215;  #10 
a = 8'd126; b = 8'd216;  #10 
a = 8'd126; b = 8'd217;  #10 
a = 8'd126; b = 8'd218;  #10 
a = 8'd126; b = 8'd219;  #10 
a = 8'd126; b = 8'd220;  #10 
a = 8'd126; b = 8'd221;  #10 
a = 8'd126; b = 8'd222;  #10 
a = 8'd126; b = 8'd223;  #10 
a = 8'd126; b = 8'd224;  #10 
a = 8'd126; b = 8'd225;  #10 
a = 8'd126; b = 8'd226;  #10 
a = 8'd126; b = 8'd227;  #10 
a = 8'd126; b = 8'd228;  #10 
a = 8'd126; b = 8'd229;  #10 
a = 8'd126; b = 8'd230;  #10 
a = 8'd126; b = 8'd231;  #10 
a = 8'd126; b = 8'd232;  #10 
a = 8'd126; b = 8'd233;  #10 
a = 8'd126; b = 8'd234;  #10 
a = 8'd126; b = 8'd235;  #10 
a = 8'd126; b = 8'd236;  #10 
a = 8'd126; b = 8'd237;  #10 
a = 8'd126; b = 8'd238;  #10 
a = 8'd126; b = 8'd239;  #10 
a = 8'd126; b = 8'd240;  #10 
a = 8'd126; b = 8'd241;  #10 
a = 8'd126; b = 8'd242;  #10 
a = 8'd126; b = 8'd243;  #10 
a = 8'd126; b = 8'd244;  #10 
a = 8'd126; b = 8'd245;  #10 
a = 8'd126; b = 8'd246;  #10 
a = 8'd126; b = 8'd247;  #10 
a = 8'd126; b = 8'd248;  #10 
a = 8'd126; b = 8'd249;  #10 
a = 8'd126; b = 8'd250;  #10 
a = 8'd126; b = 8'd251;  #10 
a = 8'd126; b = 8'd252;  #10 
a = 8'd126; b = 8'd253;  #10 
a = 8'd126; b = 8'd254;  #10 
a = 8'd126; b = 8'd255;  #10 
a = 8'd127; b = 8'd0;  #10 
a = 8'd127; b = 8'd1;  #10 
a = 8'd127; b = 8'd2;  #10 
a = 8'd127; b = 8'd3;  #10 
a = 8'd127; b = 8'd4;  #10 
a = 8'd127; b = 8'd5;  #10 
a = 8'd127; b = 8'd6;  #10 
a = 8'd127; b = 8'd7;  #10 
a = 8'd127; b = 8'd8;  #10 
a = 8'd127; b = 8'd9;  #10 
a = 8'd127; b = 8'd10;  #10 
a = 8'd127; b = 8'd11;  #10 
a = 8'd127; b = 8'd12;  #10 
a = 8'd127; b = 8'd13;  #10 
a = 8'd127; b = 8'd14;  #10 
a = 8'd127; b = 8'd15;  #10 
a = 8'd127; b = 8'd16;  #10 
a = 8'd127; b = 8'd17;  #10 
a = 8'd127; b = 8'd18;  #10 
a = 8'd127; b = 8'd19;  #10 
a = 8'd127; b = 8'd20;  #10 
a = 8'd127; b = 8'd21;  #10 
a = 8'd127; b = 8'd22;  #10 
a = 8'd127; b = 8'd23;  #10 
a = 8'd127; b = 8'd24;  #10 
a = 8'd127; b = 8'd25;  #10 
a = 8'd127; b = 8'd26;  #10 
a = 8'd127; b = 8'd27;  #10 
a = 8'd127; b = 8'd28;  #10 
a = 8'd127; b = 8'd29;  #10 
a = 8'd127; b = 8'd30;  #10 
a = 8'd127; b = 8'd31;  #10 
a = 8'd127; b = 8'd32;  #10 
a = 8'd127; b = 8'd33;  #10 
a = 8'd127; b = 8'd34;  #10 
a = 8'd127; b = 8'd35;  #10 
a = 8'd127; b = 8'd36;  #10 
a = 8'd127; b = 8'd37;  #10 
a = 8'd127; b = 8'd38;  #10 
a = 8'd127; b = 8'd39;  #10 
a = 8'd127; b = 8'd40;  #10 
a = 8'd127; b = 8'd41;  #10 
a = 8'd127; b = 8'd42;  #10 
a = 8'd127; b = 8'd43;  #10 
a = 8'd127; b = 8'd44;  #10 
a = 8'd127; b = 8'd45;  #10 
a = 8'd127; b = 8'd46;  #10 
a = 8'd127; b = 8'd47;  #10 
a = 8'd127; b = 8'd48;  #10 
a = 8'd127; b = 8'd49;  #10 
a = 8'd127; b = 8'd50;  #10 
a = 8'd127; b = 8'd51;  #10 
a = 8'd127; b = 8'd52;  #10 
a = 8'd127; b = 8'd53;  #10 
a = 8'd127; b = 8'd54;  #10 
a = 8'd127; b = 8'd55;  #10 
a = 8'd127; b = 8'd56;  #10 
a = 8'd127; b = 8'd57;  #10 
a = 8'd127; b = 8'd58;  #10 
a = 8'd127; b = 8'd59;  #10 
a = 8'd127; b = 8'd60;  #10 
a = 8'd127; b = 8'd61;  #10 
a = 8'd127; b = 8'd62;  #10 
a = 8'd127; b = 8'd63;  #10 
a = 8'd127; b = 8'd64;  #10 
a = 8'd127; b = 8'd65;  #10 
a = 8'd127; b = 8'd66;  #10 
a = 8'd127; b = 8'd67;  #10 
a = 8'd127; b = 8'd68;  #10 
a = 8'd127; b = 8'd69;  #10 
a = 8'd127; b = 8'd70;  #10 
a = 8'd127; b = 8'd71;  #10 
a = 8'd127; b = 8'd72;  #10 
a = 8'd127; b = 8'd73;  #10 
a = 8'd127; b = 8'd74;  #10 
a = 8'd127; b = 8'd75;  #10 
a = 8'd127; b = 8'd76;  #10 
a = 8'd127; b = 8'd77;  #10 
a = 8'd127; b = 8'd78;  #10 
a = 8'd127; b = 8'd79;  #10 
a = 8'd127; b = 8'd80;  #10 
a = 8'd127; b = 8'd81;  #10 
a = 8'd127; b = 8'd82;  #10 
a = 8'd127; b = 8'd83;  #10 
a = 8'd127; b = 8'd84;  #10 
a = 8'd127; b = 8'd85;  #10 
a = 8'd127; b = 8'd86;  #10 
a = 8'd127; b = 8'd87;  #10 
a = 8'd127; b = 8'd88;  #10 
a = 8'd127; b = 8'd89;  #10 
a = 8'd127; b = 8'd90;  #10 
a = 8'd127; b = 8'd91;  #10 
a = 8'd127; b = 8'd92;  #10 
a = 8'd127; b = 8'd93;  #10 
a = 8'd127; b = 8'd94;  #10 
a = 8'd127; b = 8'd95;  #10 
a = 8'd127; b = 8'd96;  #10 
a = 8'd127; b = 8'd97;  #10 
a = 8'd127; b = 8'd98;  #10 
a = 8'd127; b = 8'd99;  #10 
a = 8'd127; b = 8'd100;  #10 
a = 8'd127; b = 8'd101;  #10 
a = 8'd127; b = 8'd102;  #10 
a = 8'd127; b = 8'd103;  #10 
a = 8'd127; b = 8'd104;  #10 
a = 8'd127; b = 8'd105;  #10 
a = 8'd127; b = 8'd106;  #10 
a = 8'd127; b = 8'd107;  #10 
a = 8'd127; b = 8'd108;  #10 
a = 8'd127; b = 8'd109;  #10 
a = 8'd127; b = 8'd110;  #10 
a = 8'd127; b = 8'd111;  #10 
a = 8'd127; b = 8'd112;  #10 
a = 8'd127; b = 8'd113;  #10 
a = 8'd127; b = 8'd114;  #10 
a = 8'd127; b = 8'd115;  #10 
a = 8'd127; b = 8'd116;  #10 
a = 8'd127; b = 8'd117;  #10 
a = 8'd127; b = 8'd118;  #10 
a = 8'd127; b = 8'd119;  #10 
a = 8'd127; b = 8'd120;  #10 
a = 8'd127; b = 8'd121;  #10 
a = 8'd127; b = 8'd122;  #10 
a = 8'd127; b = 8'd123;  #10 
a = 8'd127; b = 8'd124;  #10 
a = 8'd127; b = 8'd125;  #10 
a = 8'd127; b = 8'd126;  #10 
a = 8'd127; b = 8'd127;  #10 
a = 8'd127; b = 8'd128;  #10 
a = 8'd127; b = 8'd129;  #10 
a = 8'd127; b = 8'd130;  #10 
a = 8'd127; b = 8'd131;  #10 
a = 8'd127; b = 8'd132;  #10 
a = 8'd127; b = 8'd133;  #10 
a = 8'd127; b = 8'd134;  #10 
a = 8'd127; b = 8'd135;  #10 
a = 8'd127; b = 8'd136;  #10 
a = 8'd127; b = 8'd137;  #10 
a = 8'd127; b = 8'd138;  #10 
a = 8'd127; b = 8'd139;  #10 
a = 8'd127; b = 8'd140;  #10 
a = 8'd127; b = 8'd141;  #10 
a = 8'd127; b = 8'd142;  #10 
a = 8'd127; b = 8'd143;  #10 
a = 8'd127; b = 8'd144;  #10 
a = 8'd127; b = 8'd145;  #10 
a = 8'd127; b = 8'd146;  #10 
a = 8'd127; b = 8'd147;  #10 
a = 8'd127; b = 8'd148;  #10 
a = 8'd127; b = 8'd149;  #10 
a = 8'd127; b = 8'd150;  #10 
a = 8'd127; b = 8'd151;  #10 
a = 8'd127; b = 8'd152;  #10 
a = 8'd127; b = 8'd153;  #10 
a = 8'd127; b = 8'd154;  #10 
a = 8'd127; b = 8'd155;  #10 
a = 8'd127; b = 8'd156;  #10 
a = 8'd127; b = 8'd157;  #10 
a = 8'd127; b = 8'd158;  #10 
a = 8'd127; b = 8'd159;  #10 
a = 8'd127; b = 8'd160;  #10 
a = 8'd127; b = 8'd161;  #10 
a = 8'd127; b = 8'd162;  #10 
a = 8'd127; b = 8'd163;  #10 
a = 8'd127; b = 8'd164;  #10 
a = 8'd127; b = 8'd165;  #10 
a = 8'd127; b = 8'd166;  #10 
a = 8'd127; b = 8'd167;  #10 
a = 8'd127; b = 8'd168;  #10 
a = 8'd127; b = 8'd169;  #10 
a = 8'd127; b = 8'd170;  #10 
a = 8'd127; b = 8'd171;  #10 
a = 8'd127; b = 8'd172;  #10 
a = 8'd127; b = 8'd173;  #10 
a = 8'd127; b = 8'd174;  #10 
a = 8'd127; b = 8'd175;  #10 
a = 8'd127; b = 8'd176;  #10 
a = 8'd127; b = 8'd177;  #10 
a = 8'd127; b = 8'd178;  #10 
a = 8'd127; b = 8'd179;  #10 
a = 8'd127; b = 8'd180;  #10 
a = 8'd127; b = 8'd181;  #10 
a = 8'd127; b = 8'd182;  #10 
a = 8'd127; b = 8'd183;  #10 
a = 8'd127; b = 8'd184;  #10 
a = 8'd127; b = 8'd185;  #10 
a = 8'd127; b = 8'd186;  #10 
a = 8'd127; b = 8'd187;  #10 
a = 8'd127; b = 8'd188;  #10 
a = 8'd127; b = 8'd189;  #10 
a = 8'd127; b = 8'd190;  #10 
a = 8'd127; b = 8'd191;  #10 
a = 8'd127; b = 8'd192;  #10 
a = 8'd127; b = 8'd193;  #10 
a = 8'd127; b = 8'd194;  #10 
a = 8'd127; b = 8'd195;  #10 
a = 8'd127; b = 8'd196;  #10 
a = 8'd127; b = 8'd197;  #10 
a = 8'd127; b = 8'd198;  #10 
a = 8'd127; b = 8'd199;  #10 
a = 8'd127; b = 8'd200;  #10 
a = 8'd127; b = 8'd201;  #10 
a = 8'd127; b = 8'd202;  #10 
a = 8'd127; b = 8'd203;  #10 
a = 8'd127; b = 8'd204;  #10 
a = 8'd127; b = 8'd205;  #10 
a = 8'd127; b = 8'd206;  #10 
a = 8'd127; b = 8'd207;  #10 
a = 8'd127; b = 8'd208;  #10 
a = 8'd127; b = 8'd209;  #10 
a = 8'd127; b = 8'd210;  #10 
a = 8'd127; b = 8'd211;  #10 
a = 8'd127; b = 8'd212;  #10 
a = 8'd127; b = 8'd213;  #10 
a = 8'd127; b = 8'd214;  #10 
a = 8'd127; b = 8'd215;  #10 
a = 8'd127; b = 8'd216;  #10 
a = 8'd127; b = 8'd217;  #10 
a = 8'd127; b = 8'd218;  #10 
a = 8'd127; b = 8'd219;  #10 
a = 8'd127; b = 8'd220;  #10 
a = 8'd127; b = 8'd221;  #10 
a = 8'd127; b = 8'd222;  #10 
a = 8'd127; b = 8'd223;  #10 
a = 8'd127; b = 8'd224;  #10 
a = 8'd127; b = 8'd225;  #10 
a = 8'd127; b = 8'd226;  #10 
a = 8'd127; b = 8'd227;  #10 
a = 8'd127; b = 8'd228;  #10 
a = 8'd127; b = 8'd229;  #10 
a = 8'd127; b = 8'd230;  #10 
a = 8'd127; b = 8'd231;  #10 
a = 8'd127; b = 8'd232;  #10 
a = 8'd127; b = 8'd233;  #10 
a = 8'd127; b = 8'd234;  #10 
a = 8'd127; b = 8'd235;  #10 
a = 8'd127; b = 8'd236;  #10 
a = 8'd127; b = 8'd237;  #10 
a = 8'd127; b = 8'd238;  #10 
a = 8'd127; b = 8'd239;  #10 
a = 8'd127; b = 8'd240;  #10 
a = 8'd127; b = 8'd241;  #10 
a = 8'd127; b = 8'd242;  #10 
a = 8'd127; b = 8'd243;  #10 
a = 8'd127; b = 8'd244;  #10 
a = 8'd127; b = 8'd245;  #10 
a = 8'd127; b = 8'd246;  #10 
a = 8'd127; b = 8'd247;  #10 
a = 8'd127; b = 8'd248;  #10 
a = 8'd127; b = 8'd249;  #10 
a = 8'd127; b = 8'd250;  #10 
a = 8'd127; b = 8'd251;  #10 
a = 8'd127; b = 8'd252;  #10 
a = 8'd127; b = 8'd253;  #10 
a = 8'd127; b = 8'd254;  #10 
a = 8'd127; b = 8'd255;  #10 
a = 8'd128; b = 8'd0;  #10 
a = 8'd128; b = 8'd1;  #10 
a = 8'd128; b = 8'd2;  #10 
a = 8'd128; b = 8'd3;  #10 
a = 8'd128; b = 8'd4;  #10 
a = 8'd128; b = 8'd5;  #10 
a = 8'd128; b = 8'd6;  #10 
a = 8'd128; b = 8'd7;  #10 
a = 8'd128; b = 8'd8;  #10 
a = 8'd128; b = 8'd9;  #10 
a = 8'd128; b = 8'd10;  #10 
a = 8'd128; b = 8'd11;  #10 
a = 8'd128; b = 8'd12;  #10 
a = 8'd128; b = 8'd13;  #10 
a = 8'd128; b = 8'd14;  #10 
a = 8'd128; b = 8'd15;  #10 
a = 8'd128; b = 8'd16;  #10 
a = 8'd128; b = 8'd17;  #10 
a = 8'd128; b = 8'd18;  #10 
a = 8'd128; b = 8'd19;  #10 
a = 8'd128; b = 8'd20;  #10 
a = 8'd128; b = 8'd21;  #10 
a = 8'd128; b = 8'd22;  #10 
a = 8'd128; b = 8'd23;  #10 
a = 8'd128; b = 8'd24;  #10 
a = 8'd128; b = 8'd25;  #10 
a = 8'd128; b = 8'd26;  #10 
a = 8'd128; b = 8'd27;  #10 
a = 8'd128; b = 8'd28;  #10 
a = 8'd128; b = 8'd29;  #10 
a = 8'd128; b = 8'd30;  #10 
a = 8'd128; b = 8'd31;  #10 
a = 8'd128; b = 8'd32;  #10 
a = 8'd128; b = 8'd33;  #10 
a = 8'd128; b = 8'd34;  #10 
a = 8'd128; b = 8'd35;  #10 
a = 8'd128; b = 8'd36;  #10 
a = 8'd128; b = 8'd37;  #10 
a = 8'd128; b = 8'd38;  #10 
a = 8'd128; b = 8'd39;  #10 
a = 8'd128; b = 8'd40;  #10 
a = 8'd128; b = 8'd41;  #10 
a = 8'd128; b = 8'd42;  #10 
a = 8'd128; b = 8'd43;  #10 
a = 8'd128; b = 8'd44;  #10 
a = 8'd128; b = 8'd45;  #10 
a = 8'd128; b = 8'd46;  #10 
a = 8'd128; b = 8'd47;  #10 
a = 8'd128; b = 8'd48;  #10 
a = 8'd128; b = 8'd49;  #10 
a = 8'd128; b = 8'd50;  #10 
a = 8'd128; b = 8'd51;  #10 
a = 8'd128; b = 8'd52;  #10 
a = 8'd128; b = 8'd53;  #10 
a = 8'd128; b = 8'd54;  #10 
a = 8'd128; b = 8'd55;  #10 
a = 8'd128; b = 8'd56;  #10 
a = 8'd128; b = 8'd57;  #10 
a = 8'd128; b = 8'd58;  #10 
a = 8'd128; b = 8'd59;  #10 
a = 8'd128; b = 8'd60;  #10 
a = 8'd128; b = 8'd61;  #10 
a = 8'd128; b = 8'd62;  #10 
a = 8'd128; b = 8'd63;  #10 
a = 8'd128; b = 8'd64;  #10 
a = 8'd128; b = 8'd65;  #10 
a = 8'd128; b = 8'd66;  #10 
a = 8'd128; b = 8'd67;  #10 
a = 8'd128; b = 8'd68;  #10 
a = 8'd128; b = 8'd69;  #10 
a = 8'd128; b = 8'd70;  #10 
a = 8'd128; b = 8'd71;  #10 
a = 8'd128; b = 8'd72;  #10 
a = 8'd128; b = 8'd73;  #10 
a = 8'd128; b = 8'd74;  #10 
a = 8'd128; b = 8'd75;  #10 
a = 8'd128; b = 8'd76;  #10 
a = 8'd128; b = 8'd77;  #10 
a = 8'd128; b = 8'd78;  #10 
a = 8'd128; b = 8'd79;  #10 
a = 8'd128; b = 8'd80;  #10 
a = 8'd128; b = 8'd81;  #10 
a = 8'd128; b = 8'd82;  #10 
a = 8'd128; b = 8'd83;  #10 
a = 8'd128; b = 8'd84;  #10 
a = 8'd128; b = 8'd85;  #10 
a = 8'd128; b = 8'd86;  #10 
a = 8'd128; b = 8'd87;  #10 
a = 8'd128; b = 8'd88;  #10 
a = 8'd128; b = 8'd89;  #10 
a = 8'd128; b = 8'd90;  #10 
a = 8'd128; b = 8'd91;  #10 
a = 8'd128; b = 8'd92;  #10 
a = 8'd128; b = 8'd93;  #10 
a = 8'd128; b = 8'd94;  #10 
a = 8'd128; b = 8'd95;  #10 
a = 8'd128; b = 8'd96;  #10 
a = 8'd128; b = 8'd97;  #10 
a = 8'd128; b = 8'd98;  #10 
a = 8'd128; b = 8'd99;  #10 
a = 8'd128; b = 8'd100;  #10 
a = 8'd128; b = 8'd101;  #10 
a = 8'd128; b = 8'd102;  #10 
a = 8'd128; b = 8'd103;  #10 
a = 8'd128; b = 8'd104;  #10 
a = 8'd128; b = 8'd105;  #10 
a = 8'd128; b = 8'd106;  #10 
a = 8'd128; b = 8'd107;  #10 
a = 8'd128; b = 8'd108;  #10 
a = 8'd128; b = 8'd109;  #10 
a = 8'd128; b = 8'd110;  #10 
a = 8'd128; b = 8'd111;  #10 
a = 8'd128; b = 8'd112;  #10 
a = 8'd128; b = 8'd113;  #10 
a = 8'd128; b = 8'd114;  #10 
a = 8'd128; b = 8'd115;  #10 
a = 8'd128; b = 8'd116;  #10 
a = 8'd128; b = 8'd117;  #10 
a = 8'd128; b = 8'd118;  #10 
a = 8'd128; b = 8'd119;  #10 
a = 8'd128; b = 8'd120;  #10 
a = 8'd128; b = 8'd121;  #10 
a = 8'd128; b = 8'd122;  #10 
a = 8'd128; b = 8'd123;  #10 
a = 8'd128; b = 8'd124;  #10 
a = 8'd128; b = 8'd125;  #10 
a = 8'd128; b = 8'd126;  #10 
a = 8'd128; b = 8'd127;  #10 
a = 8'd128; b = 8'd128;  #10 
a = 8'd128; b = 8'd129;  #10 
a = 8'd128; b = 8'd130;  #10 
a = 8'd128; b = 8'd131;  #10 
a = 8'd128; b = 8'd132;  #10 
a = 8'd128; b = 8'd133;  #10 
a = 8'd128; b = 8'd134;  #10 
a = 8'd128; b = 8'd135;  #10 
a = 8'd128; b = 8'd136;  #10 
a = 8'd128; b = 8'd137;  #10 
a = 8'd128; b = 8'd138;  #10 
a = 8'd128; b = 8'd139;  #10 
a = 8'd128; b = 8'd140;  #10 
a = 8'd128; b = 8'd141;  #10 
a = 8'd128; b = 8'd142;  #10 
a = 8'd128; b = 8'd143;  #10 
a = 8'd128; b = 8'd144;  #10 
a = 8'd128; b = 8'd145;  #10 
a = 8'd128; b = 8'd146;  #10 
a = 8'd128; b = 8'd147;  #10 
a = 8'd128; b = 8'd148;  #10 
a = 8'd128; b = 8'd149;  #10 
a = 8'd128; b = 8'd150;  #10 
a = 8'd128; b = 8'd151;  #10 
a = 8'd128; b = 8'd152;  #10 
a = 8'd128; b = 8'd153;  #10 
a = 8'd128; b = 8'd154;  #10 
a = 8'd128; b = 8'd155;  #10 
a = 8'd128; b = 8'd156;  #10 
a = 8'd128; b = 8'd157;  #10 
a = 8'd128; b = 8'd158;  #10 
a = 8'd128; b = 8'd159;  #10 
a = 8'd128; b = 8'd160;  #10 
a = 8'd128; b = 8'd161;  #10 
a = 8'd128; b = 8'd162;  #10 
a = 8'd128; b = 8'd163;  #10 
a = 8'd128; b = 8'd164;  #10 
a = 8'd128; b = 8'd165;  #10 
a = 8'd128; b = 8'd166;  #10 
a = 8'd128; b = 8'd167;  #10 
a = 8'd128; b = 8'd168;  #10 
a = 8'd128; b = 8'd169;  #10 
a = 8'd128; b = 8'd170;  #10 
a = 8'd128; b = 8'd171;  #10 
a = 8'd128; b = 8'd172;  #10 
a = 8'd128; b = 8'd173;  #10 
a = 8'd128; b = 8'd174;  #10 
a = 8'd128; b = 8'd175;  #10 
a = 8'd128; b = 8'd176;  #10 
a = 8'd128; b = 8'd177;  #10 
a = 8'd128; b = 8'd178;  #10 
a = 8'd128; b = 8'd179;  #10 
a = 8'd128; b = 8'd180;  #10 
a = 8'd128; b = 8'd181;  #10 
a = 8'd128; b = 8'd182;  #10 
a = 8'd128; b = 8'd183;  #10 
a = 8'd128; b = 8'd184;  #10 
a = 8'd128; b = 8'd185;  #10 
a = 8'd128; b = 8'd186;  #10 
a = 8'd128; b = 8'd187;  #10 
a = 8'd128; b = 8'd188;  #10 
a = 8'd128; b = 8'd189;  #10 
a = 8'd128; b = 8'd190;  #10 
a = 8'd128; b = 8'd191;  #10 
a = 8'd128; b = 8'd192;  #10 
a = 8'd128; b = 8'd193;  #10 
a = 8'd128; b = 8'd194;  #10 
a = 8'd128; b = 8'd195;  #10 
a = 8'd128; b = 8'd196;  #10 
a = 8'd128; b = 8'd197;  #10 
a = 8'd128; b = 8'd198;  #10 
a = 8'd128; b = 8'd199;  #10 
a = 8'd128; b = 8'd200;  #10 
a = 8'd128; b = 8'd201;  #10 
a = 8'd128; b = 8'd202;  #10 
a = 8'd128; b = 8'd203;  #10 
a = 8'd128; b = 8'd204;  #10 
a = 8'd128; b = 8'd205;  #10 
a = 8'd128; b = 8'd206;  #10 
a = 8'd128; b = 8'd207;  #10 
a = 8'd128; b = 8'd208;  #10 
a = 8'd128; b = 8'd209;  #10 
a = 8'd128; b = 8'd210;  #10 
a = 8'd128; b = 8'd211;  #10 
a = 8'd128; b = 8'd212;  #10 
a = 8'd128; b = 8'd213;  #10 
a = 8'd128; b = 8'd214;  #10 
a = 8'd128; b = 8'd215;  #10 
a = 8'd128; b = 8'd216;  #10 
a = 8'd128; b = 8'd217;  #10 
a = 8'd128; b = 8'd218;  #10 
a = 8'd128; b = 8'd219;  #10 
a = 8'd128; b = 8'd220;  #10 
a = 8'd128; b = 8'd221;  #10 
a = 8'd128; b = 8'd222;  #10 
a = 8'd128; b = 8'd223;  #10 
a = 8'd128; b = 8'd224;  #10 
a = 8'd128; b = 8'd225;  #10 
a = 8'd128; b = 8'd226;  #10 
a = 8'd128; b = 8'd227;  #10 
a = 8'd128; b = 8'd228;  #10 
a = 8'd128; b = 8'd229;  #10 
a = 8'd128; b = 8'd230;  #10 
a = 8'd128; b = 8'd231;  #10 
a = 8'd128; b = 8'd232;  #10 
a = 8'd128; b = 8'd233;  #10 
a = 8'd128; b = 8'd234;  #10 
a = 8'd128; b = 8'd235;  #10 
a = 8'd128; b = 8'd236;  #10 
a = 8'd128; b = 8'd237;  #10 
a = 8'd128; b = 8'd238;  #10 
a = 8'd128; b = 8'd239;  #10 
a = 8'd128; b = 8'd240;  #10 
a = 8'd128; b = 8'd241;  #10 
a = 8'd128; b = 8'd242;  #10 
a = 8'd128; b = 8'd243;  #10 
a = 8'd128; b = 8'd244;  #10 
a = 8'd128; b = 8'd245;  #10 
a = 8'd128; b = 8'd246;  #10 
a = 8'd128; b = 8'd247;  #10 
a = 8'd128; b = 8'd248;  #10 
a = 8'd128; b = 8'd249;  #10 
a = 8'd128; b = 8'd250;  #10 
a = 8'd128; b = 8'd251;  #10 
a = 8'd128; b = 8'd252;  #10 
a = 8'd128; b = 8'd253;  #10 
a = 8'd128; b = 8'd254;  #10 
a = 8'd128; b = 8'd255;  #10 
a = 8'd129; b = 8'd0;  #10 
a = 8'd129; b = 8'd1;  #10 
a = 8'd129; b = 8'd2;  #10 
a = 8'd129; b = 8'd3;  #10 
a = 8'd129; b = 8'd4;  #10 
a = 8'd129; b = 8'd5;  #10 
a = 8'd129; b = 8'd6;  #10 
a = 8'd129; b = 8'd7;  #10 
a = 8'd129; b = 8'd8;  #10 
a = 8'd129; b = 8'd9;  #10 
a = 8'd129; b = 8'd10;  #10 
a = 8'd129; b = 8'd11;  #10 
a = 8'd129; b = 8'd12;  #10 
a = 8'd129; b = 8'd13;  #10 
a = 8'd129; b = 8'd14;  #10 
a = 8'd129; b = 8'd15;  #10 
a = 8'd129; b = 8'd16;  #10 
a = 8'd129; b = 8'd17;  #10 
a = 8'd129; b = 8'd18;  #10 
a = 8'd129; b = 8'd19;  #10 
a = 8'd129; b = 8'd20;  #10 
a = 8'd129; b = 8'd21;  #10 
a = 8'd129; b = 8'd22;  #10 
a = 8'd129; b = 8'd23;  #10 
a = 8'd129; b = 8'd24;  #10 
a = 8'd129; b = 8'd25;  #10 
a = 8'd129; b = 8'd26;  #10 
a = 8'd129; b = 8'd27;  #10 
a = 8'd129; b = 8'd28;  #10 
a = 8'd129; b = 8'd29;  #10 
a = 8'd129; b = 8'd30;  #10 
a = 8'd129; b = 8'd31;  #10 
a = 8'd129; b = 8'd32;  #10 
a = 8'd129; b = 8'd33;  #10 
a = 8'd129; b = 8'd34;  #10 
a = 8'd129; b = 8'd35;  #10 
a = 8'd129; b = 8'd36;  #10 
a = 8'd129; b = 8'd37;  #10 
a = 8'd129; b = 8'd38;  #10 
a = 8'd129; b = 8'd39;  #10 
a = 8'd129; b = 8'd40;  #10 
a = 8'd129; b = 8'd41;  #10 
a = 8'd129; b = 8'd42;  #10 
a = 8'd129; b = 8'd43;  #10 
a = 8'd129; b = 8'd44;  #10 
a = 8'd129; b = 8'd45;  #10 
a = 8'd129; b = 8'd46;  #10 
a = 8'd129; b = 8'd47;  #10 
a = 8'd129; b = 8'd48;  #10 
a = 8'd129; b = 8'd49;  #10 
a = 8'd129; b = 8'd50;  #10 
a = 8'd129; b = 8'd51;  #10 
a = 8'd129; b = 8'd52;  #10 
a = 8'd129; b = 8'd53;  #10 
a = 8'd129; b = 8'd54;  #10 
a = 8'd129; b = 8'd55;  #10 
a = 8'd129; b = 8'd56;  #10 
a = 8'd129; b = 8'd57;  #10 
a = 8'd129; b = 8'd58;  #10 
a = 8'd129; b = 8'd59;  #10 
a = 8'd129; b = 8'd60;  #10 
a = 8'd129; b = 8'd61;  #10 
a = 8'd129; b = 8'd62;  #10 
a = 8'd129; b = 8'd63;  #10 
a = 8'd129; b = 8'd64;  #10 
a = 8'd129; b = 8'd65;  #10 
a = 8'd129; b = 8'd66;  #10 
a = 8'd129; b = 8'd67;  #10 
a = 8'd129; b = 8'd68;  #10 
a = 8'd129; b = 8'd69;  #10 
a = 8'd129; b = 8'd70;  #10 
a = 8'd129; b = 8'd71;  #10 
a = 8'd129; b = 8'd72;  #10 
a = 8'd129; b = 8'd73;  #10 
a = 8'd129; b = 8'd74;  #10 
a = 8'd129; b = 8'd75;  #10 
a = 8'd129; b = 8'd76;  #10 
a = 8'd129; b = 8'd77;  #10 
a = 8'd129; b = 8'd78;  #10 
a = 8'd129; b = 8'd79;  #10 
a = 8'd129; b = 8'd80;  #10 
a = 8'd129; b = 8'd81;  #10 
a = 8'd129; b = 8'd82;  #10 
a = 8'd129; b = 8'd83;  #10 
a = 8'd129; b = 8'd84;  #10 
a = 8'd129; b = 8'd85;  #10 
a = 8'd129; b = 8'd86;  #10 
a = 8'd129; b = 8'd87;  #10 
a = 8'd129; b = 8'd88;  #10 
a = 8'd129; b = 8'd89;  #10 
a = 8'd129; b = 8'd90;  #10 
a = 8'd129; b = 8'd91;  #10 
a = 8'd129; b = 8'd92;  #10 
a = 8'd129; b = 8'd93;  #10 
a = 8'd129; b = 8'd94;  #10 
a = 8'd129; b = 8'd95;  #10 
a = 8'd129; b = 8'd96;  #10 
a = 8'd129; b = 8'd97;  #10 
a = 8'd129; b = 8'd98;  #10 
a = 8'd129; b = 8'd99;  #10 
a = 8'd129; b = 8'd100;  #10 
a = 8'd129; b = 8'd101;  #10 
a = 8'd129; b = 8'd102;  #10 
a = 8'd129; b = 8'd103;  #10 
a = 8'd129; b = 8'd104;  #10 
a = 8'd129; b = 8'd105;  #10 
a = 8'd129; b = 8'd106;  #10 
a = 8'd129; b = 8'd107;  #10 
a = 8'd129; b = 8'd108;  #10 
a = 8'd129; b = 8'd109;  #10 
a = 8'd129; b = 8'd110;  #10 
a = 8'd129; b = 8'd111;  #10 
a = 8'd129; b = 8'd112;  #10 
a = 8'd129; b = 8'd113;  #10 
a = 8'd129; b = 8'd114;  #10 
a = 8'd129; b = 8'd115;  #10 
a = 8'd129; b = 8'd116;  #10 
a = 8'd129; b = 8'd117;  #10 
a = 8'd129; b = 8'd118;  #10 
a = 8'd129; b = 8'd119;  #10 
a = 8'd129; b = 8'd120;  #10 
a = 8'd129; b = 8'd121;  #10 
a = 8'd129; b = 8'd122;  #10 
a = 8'd129; b = 8'd123;  #10 
a = 8'd129; b = 8'd124;  #10 
a = 8'd129; b = 8'd125;  #10 
a = 8'd129; b = 8'd126;  #10 
a = 8'd129; b = 8'd127;  #10 
a = 8'd129; b = 8'd128;  #10 
a = 8'd129; b = 8'd129;  #10 
a = 8'd129; b = 8'd130;  #10 
a = 8'd129; b = 8'd131;  #10 
a = 8'd129; b = 8'd132;  #10 
a = 8'd129; b = 8'd133;  #10 
a = 8'd129; b = 8'd134;  #10 
a = 8'd129; b = 8'd135;  #10 
a = 8'd129; b = 8'd136;  #10 
a = 8'd129; b = 8'd137;  #10 
a = 8'd129; b = 8'd138;  #10 
a = 8'd129; b = 8'd139;  #10 
a = 8'd129; b = 8'd140;  #10 
a = 8'd129; b = 8'd141;  #10 
a = 8'd129; b = 8'd142;  #10 
a = 8'd129; b = 8'd143;  #10 
a = 8'd129; b = 8'd144;  #10 
a = 8'd129; b = 8'd145;  #10 
a = 8'd129; b = 8'd146;  #10 
a = 8'd129; b = 8'd147;  #10 
a = 8'd129; b = 8'd148;  #10 
a = 8'd129; b = 8'd149;  #10 
a = 8'd129; b = 8'd150;  #10 
a = 8'd129; b = 8'd151;  #10 
a = 8'd129; b = 8'd152;  #10 
a = 8'd129; b = 8'd153;  #10 
a = 8'd129; b = 8'd154;  #10 
a = 8'd129; b = 8'd155;  #10 
a = 8'd129; b = 8'd156;  #10 
a = 8'd129; b = 8'd157;  #10 
a = 8'd129; b = 8'd158;  #10 
a = 8'd129; b = 8'd159;  #10 
a = 8'd129; b = 8'd160;  #10 
a = 8'd129; b = 8'd161;  #10 
a = 8'd129; b = 8'd162;  #10 
a = 8'd129; b = 8'd163;  #10 
a = 8'd129; b = 8'd164;  #10 
a = 8'd129; b = 8'd165;  #10 
a = 8'd129; b = 8'd166;  #10 
a = 8'd129; b = 8'd167;  #10 
a = 8'd129; b = 8'd168;  #10 
a = 8'd129; b = 8'd169;  #10 
a = 8'd129; b = 8'd170;  #10 
a = 8'd129; b = 8'd171;  #10 
a = 8'd129; b = 8'd172;  #10 
a = 8'd129; b = 8'd173;  #10 
a = 8'd129; b = 8'd174;  #10 
a = 8'd129; b = 8'd175;  #10 
a = 8'd129; b = 8'd176;  #10 
a = 8'd129; b = 8'd177;  #10 
a = 8'd129; b = 8'd178;  #10 
a = 8'd129; b = 8'd179;  #10 
a = 8'd129; b = 8'd180;  #10 
a = 8'd129; b = 8'd181;  #10 
a = 8'd129; b = 8'd182;  #10 
a = 8'd129; b = 8'd183;  #10 
a = 8'd129; b = 8'd184;  #10 
a = 8'd129; b = 8'd185;  #10 
a = 8'd129; b = 8'd186;  #10 
a = 8'd129; b = 8'd187;  #10 
a = 8'd129; b = 8'd188;  #10 
a = 8'd129; b = 8'd189;  #10 
a = 8'd129; b = 8'd190;  #10 
a = 8'd129; b = 8'd191;  #10 
a = 8'd129; b = 8'd192;  #10 
a = 8'd129; b = 8'd193;  #10 
a = 8'd129; b = 8'd194;  #10 
a = 8'd129; b = 8'd195;  #10 
a = 8'd129; b = 8'd196;  #10 
a = 8'd129; b = 8'd197;  #10 
a = 8'd129; b = 8'd198;  #10 
a = 8'd129; b = 8'd199;  #10 
a = 8'd129; b = 8'd200;  #10 
a = 8'd129; b = 8'd201;  #10 
a = 8'd129; b = 8'd202;  #10 
a = 8'd129; b = 8'd203;  #10 
a = 8'd129; b = 8'd204;  #10 
a = 8'd129; b = 8'd205;  #10 
a = 8'd129; b = 8'd206;  #10 
a = 8'd129; b = 8'd207;  #10 
a = 8'd129; b = 8'd208;  #10 
a = 8'd129; b = 8'd209;  #10 
a = 8'd129; b = 8'd210;  #10 
a = 8'd129; b = 8'd211;  #10 
a = 8'd129; b = 8'd212;  #10 
a = 8'd129; b = 8'd213;  #10 
a = 8'd129; b = 8'd214;  #10 
a = 8'd129; b = 8'd215;  #10 
a = 8'd129; b = 8'd216;  #10 
a = 8'd129; b = 8'd217;  #10 
a = 8'd129; b = 8'd218;  #10 
a = 8'd129; b = 8'd219;  #10 
a = 8'd129; b = 8'd220;  #10 
a = 8'd129; b = 8'd221;  #10 
a = 8'd129; b = 8'd222;  #10 
a = 8'd129; b = 8'd223;  #10 
a = 8'd129; b = 8'd224;  #10 
a = 8'd129; b = 8'd225;  #10 
a = 8'd129; b = 8'd226;  #10 
a = 8'd129; b = 8'd227;  #10 
a = 8'd129; b = 8'd228;  #10 
a = 8'd129; b = 8'd229;  #10 
a = 8'd129; b = 8'd230;  #10 
a = 8'd129; b = 8'd231;  #10 
a = 8'd129; b = 8'd232;  #10 
a = 8'd129; b = 8'd233;  #10 
a = 8'd129; b = 8'd234;  #10 
a = 8'd129; b = 8'd235;  #10 
a = 8'd129; b = 8'd236;  #10 
a = 8'd129; b = 8'd237;  #10 
a = 8'd129; b = 8'd238;  #10 
a = 8'd129; b = 8'd239;  #10 
a = 8'd129; b = 8'd240;  #10 
a = 8'd129; b = 8'd241;  #10 
a = 8'd129; b = 8'd242;  #10 
a = 8'd129; b = 8'd243;  #10 
a = 8'd129; b = 8'd244;  #10 
a = 8'd129; b = 8'd245;  #10 
a = 8'd129; b = 8'd246;  #10 
a = 8'd129; b = 8'd247;  #10 
a = 8'd129; b = 8'd248;  #10 
a = 8'd129; b = 8'd249;  #10 
a = 8'd129; b = 8'd250;  #10 
a = 8'd129; b = 8'd251;  #10 
a = 8'd129; b = 8'd252;  #10 
a = 8'd129; b = 8'd253;  #10 
a = 8'd129; b = 8'd254;  #10 
a = 8'd129; b = 8'd255;  #10 
a = 8'd130; b = 8'd0;  #10 
a = 8'd130; b = 8'd1;  #10 
a = 8'd130; b = 8'd2;  #10 
a = 8'd130; b = 8'd3;  #10 
a = 8'd130; b = 8'd4;  #10 
a = 8'd130; b = 8'd5;  #10 
a = 8'd130; b = 8'd6;  #10 
a = 8'd130; b = 8'd7;  #10 
a = 8'd130; b = 8'd8;  #10 
a = 8'd130; b = 8'd9;  #10 
a = 8'd130; b = 8'd10;  #10 
a = 8'd130; b = 8'd11;  #10 
a = 8'd130; b = 8'd12;  #10 
a = 8'd130; b = 8'd13;  #10 
a = 8'd130; b = 8'd14;  #10 
a = 8'd130; b = 8'd15;  #10 
a = 8'd130; b = 8'd16;  #10 
a = 8'd130; b = 8'd17;  #10 
a = 8'd130; b = 8'd18;  #10 
a = 8'd130; b = 8'd19;  #10 
a = 8'd130; b = 8'd20;  #10 
a = 8'd130; b = 8'd21;  #10 
a = 8'd130; b = 8'd22;  #10 
a = 8'd130; b = 8'd23;  #10 
a = 8'd130; b = 8'd24;  #10 
a = 8'd130; b = 8'd25;  #10 
a = 8'd130; b = 8'd26;  #10 
a = 8'd130; b = 8'd27;  #10 
a = 8'd130; b = 8'd28;  #10 
a = 8'd130; b = 8'd29;  #10 
a = 8'd130; b = 8'd30;  #10 
a = 8'd130; b = 8'd31;  #10 
a = 8'd130; b = 8'd32;  #10 
a = 8'd130; b = 8'd33;  #10 
a = 8'd130; b = 8'd34;  #10 
a = 8'd130; b = 8'd35;  #10 
a = 8'd130; b = 8'd36;  #10 
a = 8'd130; b = 8'd37;  #10 
a = 8'd130; b = 8'd38;  #10 
a = 8'd130; b = 8'd39;  #10 
a = 8'd130; b = 8'd40;  #10 
a = 8'd130; b = 8'd41;  #10 
a = 8'd130; b = 8'd42;  #10 
a = 8'd130; b = 8'd43;  #10 
a = 8'd130; b = 8'd44;  #10 
a = 8'd130; b = 8'd45;  #10 
a = 8'd130; b = 8'd46;  #10 
a = 8'd130; b = 8'd47;  #10 
a = 8'd130; b = 8'd48;  #10 
a = 8'd130; b = 8'd49;  #10 
a = 8'd130; b = 8'd50;  #10 
a = 8'd130; b = 8'd51;  #10 
a = 8'd130; b = 8'd52;  #10 
a = 8'd130; b = 8'd53;  #10 
a = 8'd130; b = 8'd54;  #10 
a = 8'd130; b = 8'd55;  #10 
a = 8'd130; b = 8'd56;  #10 
a = 8'd130; b = 8'd57;  #10 
a = 8'd130; b = 8'd58;  #10 
a = 8'd130; b = 8'd59;  #10 
a = 8'd130; b = 8'd60;  #10 
a = 8'd130; b = 8'd61;  #10 
a = 8'd130; b = 8'd62;  #10 
a = 8'd130; b = 8'd63;  #10 
a = 8'd130; b = 8'd64;  #10 
a = 8'd130; b = 8'd65;  #10 
a = 8'd130; b = 8'd66;  #10 
a = 8'd130; b = 8'd67;  #10 
a = 8'd130; b = 8'd68;  #10 
a = 8'd130; b = 8'd69;  #10 
a = 8'd130; b = 8'd70;  #10 
a = 8'd130; b = 8'd71;  #10 
a = 8'd130; b = 8'd72;  #10 
a = 8'd130; b = 8'd73;  #10 
a = 8'd130; b = 8'd74;  #10 
a = 8'd130; b = 8'd75;  #10 
a = 8'd130; b = 8'd76;  #10 
a = 8'd130; b = 8'd77;  #10 
a = 8'd130; b = 8'd78;  #10 
a = 8'd130; b = 8'd79;  #10 
a = 8'd130; b = 8'd80;  #10 
a = 8'd130; b = 8'd81;  #10 
a = 8'd130; b = 8'd82;  #10 
a = 8'd130; b = 8'd83;  #10 
a = 8'd130; b = 8'd84;  #10 
a = 8'd130; b = 8'd85;  #10 
a = 8'd130; b = 8'd86;  #10 
a = 8'd130; b = 8'd87;  #10 
a = 8'd130; b = 8'd88;  #10 
a = 8'd130; b = 8'd89;  #10 
a = 8'd130; b = 8'd90;  #10 
a = 8'd130; b = 8'd91;  #10 
a = 8'd130; b = 8'd92;  #10 
a = 8'd130; b = 8'd93;  #10 
a = 8'd130; b = 8'd94;  #10 
a = 8'd130; b = 8'd95;  #10 
a = 8'd130; b = 8'd96;  #10 
a = 8'd130; b = 8'd97;  #10 
a = 8'd130; b = 8'd98;  #10 
a = 8'd130; b = 8'd99;  #10 
a = 8'd130; b = 8'd100;  #10 
a = 8'd130; b = 8'd101;  #10 
a = 8'd130; b = 8'd102;  #10 
a = 8'd130; b = 8'd103;  #10 
a = 8'd130; b = 8'd104;  #10 
a = 8'd130; b = 8'd105;  #10 
a = 8'd130; b = 8'd106;  #10 
a = 8'd130; b = 8'd107;  #10 
a = 8'd130; b = 8'd108;  #10 
a = 8'd130; b = 8'd109;  #10 
a = 8'd130; b = 8'd110;  #10 
a = 8'd130; b = 8'd111;  #10 
a = 8'd130; b = 8'd112;  #10 
a = 8'd130; b = 8'd113;  #10 
a = 8'd130; b = 8'd114;  #10 
a = 8'd130; b = 8'd115;  #10 
a = 8'd130; b = 8'd116;  #10 
a = 8'd130; b = 8'd117;  #10 
a = 8'd130; b = 8'd118;  #10 
a = 8'd130; b = 8'd119;  #10 
a = 8'd130; b = 8'd120;  #10 
a = 8'd130; b = 8'd121;  #10 
a = 8'd130; b = 8'd122;  #10 
a = 8'd130; b = 8'd123;  #10 
a = 8'd130; b = 8'd124;  #10 
a = 8'd130; b = 8'd125;  #10 
a = 8'd130; b = 8'd126;  #10 
a = 8'd130; b = 8'd127;  #10 
a = 8'd130; b = 8'd128;  #10 
a = 8'd130; b = 8'd129;  #10 
a = 8'd130; b = 8'd130;  #10 
a = 8'd130; b = 8'd131;  #10 
a = 8'd130; b = 8'd132;  #10 
a = 8'd130; b = 8'd133;  #10 
a = 8'd130; b = 8'd134;  #10 
a = 8'd130; b = 8'd135;  #10 
a = 8'd130; b = 8'd136;  #10 
a = 8'd130; b = 8'd137;  #10 
a = 8'd130; b = 8'd138;  #10 
a = 8'd130; b = 8'd139;  #10 
a = 8'd130; b = 8'd140;  #10 
a = 8'd130; b = 8'd141;  #10 
a = 8'd130; b = 8'd142;  #10 
a = 8'd130; b = 8'd143;  #10 
a = 8'd130; b = 8'd144;  #10 
a = 8'd130; b = 8'd145;  #10 
a = 8'd130; b = 8'd146;  #10 
a = 8'd130; b = 8'd147;  #10 
a = 8'd130; b = 8'd148;  #10 
a = 8'd130; b = 8'd149;  #10 
a = 8'd130; b = 8'd150;  #10 
a = 8'd130; b = 8'd151;  #10 
a = 8'd130; b = 8'd152;  #10 
a = 8'd130; b = 8'd153;  #10 
a = 8'd130; b = 8'd154;  #10 
a = 8'd130; b = 8'd155;  #10 
a = 8'd130; b = 8'd156;  #10 
a = 8'd130; b = 8'd157;  #10 
a = 8'd130; b = 8'd158;  #10 
a = 8'd130; b = 8'd159;  #10 
a = 8'd130; b = 8'd160;  #10 
a = 8'd130; b = 8'd161;  #10 
a = 8'd130; b = 8'd162;  #10 
a = 8'd130; b = 8'd163;  #10 
a = 8'd130; b = 8'd164;  #10 
a = 8'd130; b = 8'd165;  #10 
a = 8'd130; b = 8'd166;  #10 
a = 8'd130; b = 8'd167;  #10 
a = 8'd130; b = 8'd168;  #10 
a = 8'd130; b = 8'd169;  #10 
a = 8'd130; b = 8'd170;  #10 
a = 8'd130; b = 8'd171;  #10 
a = 8'd130; b = 8'd172;  #10 
a = 8'd130; b = 8'd173;  #10 
a = 8'd130; b = 8'd174;  #10 
a = 8'd130; b = 8'd175;  #10 
a = 8'd130; b = 8'd176;  #10 
a = 8'd130; b = 8'd177;  #10 
a = 8'd130; b = 8'd178;  #10 
a = 8'd130; b = 8'd179;  #10 
a = 8'd130; b = 8'd180;  #10 
a = 8'd130; b = 8'd181;  #10 
a = 8'd130; b = 8'd182;  #10 
a = 8'd130; b = 8'd183;  #10 
a = 8'd130; b = 8'd184;  #10 
a = 8'd130; b = 8'd185;  #10 
a = 8'd130; b = 8'd186;  #10 
a = 8'd130; b = 8'd187;  #10 
a = 8'd130; b = 8'd188;  #10 
a = 8'd130; b = 8'd189;  #10 
a = 8'd130; b = 8'd190;  #10 
a = 8'd130; b = 8'd191;  #10 
a = 8'd130; b = 8'd192;  #10 
a = 8'd130; b = 8'd193;  #10 
a = 8'd130; b = 8'd194;  #10 
a = 8'd130; b = 8'd195;  #10 
a = 8'd130; b = 8'd196;  #10 
a = 8'd130; b = 8'd197;  #10 
a = 8'd130; b = 8'd198;  #10 
a = 8'd130; b = 8'd199;  #10 
a = 8'd130; b = 8'd200;  #10 
a = 8'd130; b = 8'd201;  #10 
a = 8'd130; b = 8'd202;  #10 
a = 8'd130; b = 8'd203;  #10 
a = 8'd130; b = 8'd204;  #10 
a = 8'd130; b = 8'd205;  #10 
a = 8'd130; b = 8'd206;  #10 
a = 8'd130; b = 8'd207;  #10 
a = 8'd130; b = 8'd208;  #10 
a = 8'd130; b = 8'd209;  #10 
a = 8'd130; b = 8'd210;  #10 
a = 8'd130; b = 8'd211;  #10 
a = 8'd130; b = 8'd212;  #10 
a = 8'd130; b = 8'd213;  #10 
a = 8'd130; b = 8'd214;  #10 
a = 8'd130; b = 8'd215;  #10 
a = 8'd130; b = 8'd216;  #10 
a = 8'd130; b = 8'd217;  #10 
a = 8'd130; b = 8'd218;  #10 
a = 8'd130; b = 8'd219;  #10 
a = 8'd130; b = 8'd220;  #10 
a = 8'd130; b = 8'd221;  #10 
a = 8'd130; b = 8'd222;  #10 
a = 8'd130; b = 8'd223;  #10 
a = 8'd130; b = 8'd224;  #10 
a = 8'd130; b = 8'd225;  #10 
a = 8'd130; b = 8'd226;  #10 
a = 8'd130; b = 8'd227;  #10 
a = 8'd130; b = 8'd228;  #10 
a = 8'd130; b = 8'd229;  #10 
a = 8'd130; b = 8'd230;  #10 
a = 8'd130; b = 8'd231;  #10 
a = 8'd130; b = 8'd232;  #10 
a = 8'd130; b = 8'd233;  #10 
a = 8'd130; b = 8'd234;  #10 
a = 8'd130; b = 8'd235;  #10 
a = 8'd130; b = 8'd236;  #10 
a = 8'd130; b = 8'd237;  #10 
a = 8'd130; b = 8'd238;  #10 
a = 8'd130; b = 8'd239;  #10 
a = 8'd130; b = 8'd240;  #10 
a = 8'd130; b = 8'd241;  #10 
a = 8'd130; b = 8'd242;  #10 
a = 8'd130; b = 8'd243;  #10 
a = 8'd130; b = 8'd244;  #10 
a = 8'd130; b = 8'd245;  #10 
a = 8'd130; b = 8'd246;  #10 
a = 8'd130; b = 8'd247;  #10 
a = 8'd130; b = 8'd248;  #10 
a = 8'd130; b = 8'd249;  #10 
a = 8'd130; b = 8'd250;  #10 
a = 8'd130; b = 8'd251;  #10 
a = 8'd130; b = 8'd252;  #10 
a = 8'd130; b = 8'd253;  #10 
a = 8'd130; b = 8'd254;  #10 
a = 8'd130; b = 8'd255;  #10 
a = 8'd131; b = 8'd0;  #10 
a = 8'd131; b = 8'd1;  #10 
a = 8'd131; b = 8'd2;  #10 
a = 8'd131; b = 8'd3;  #10 
a = 8'd131; b = 8'd4;  #10 
a = 8'd131; b = 8'd5;  #10 
a = 8'd131; b = 8'd6;  #10 
a = 8'd131; b = 8'd7;  #10 
a = 8'd131; b = 8'd8;  #10 
a = 8'd131; b = 8'd9;  #10 
a = 8'd131; b = 8'd10;  #10 
a = 8'd131; b = 8'd11;  #10 
a = 8'd131; b = 8'd12;  #10 
a = 8'd131; b = 8'd13;  #10 
a = 8'd131; b = 8'd14;  #10 
a = 8'd131; b = 8'd15;  #10 
a = 8'd131; b = 8'd16;  #10 
a = 8'd131; b = 8'd17;  #10 
a = 8'd131; b = 8'd18;  #10 
a = 8'd131; b = 8'd19;  #10 
a = 8'd131; b = 8'd20;  #10 
a = 8'd131; b = 8'd21;  #10 
a = 8'd131; b = 8'd22;  #10 
a = 8'd131; b = 8'd23;  #10 
a = 8'd131; b = 8'd24;  #10 
a = 8'd131; b = 8'd25;  #10 
a = 8'd131; b = 8'd26;  #10 
a = 8'd131; b = 8'd27;  #10 
a = 8'd131; b = 8'd28;  #10 
a = 8'd131; b = 8'd29;  #10 
a = 8'd131; b = 8'd30;  #10 
a = 8'd131; b = 8'd31;  #10 
a = 8'd131; b = 8'd32;  #10 
a = 8'd131; b = 8'd33;  #10 
a = 8'd131; b = 8'd34;  #10 
a = 8'd131; b = 8'd35;  #10 
a = 8'd131; b = 8'd36;  #10 
a = 8'd131; b = 8'd37;  #10 
a = 8'd131; b = 8'd38;  #10 
a = 8'd131; b = 8'd39;  #10 
a = 8'd131; b = 8'd40;  #10 
a = 8'd131; b = 8'd41;  #10 
a = 8'd131; b = 8'd42;  #10 
a = 8'd131; b = 8'd43;  #10 
a = 8'd131; b = 8'd44;  #10 
a = 8'd131; b = 8'd45;  #10 
a = 8'd131; b = 8'd46;  #10 
a = 8'd131; b = 8'd47;  #10 
a = 8'd131; b = 8'd48;  #10 
a = 8'd131; b = 8'd49;  #10 
a = 8'd131; b = 8'd50;  #10 
a = 8'd131; b = 8'd51;  #10 
a = 8'd131; b = 8'd52;  #10 
a = 8'd131; b = 8'd53;  #10 
a = 8'd131; b = 8'd54;  #10 
a = 8'd131; b = 8'd55;  #10 
a = 8'd131; b = 8'd56;  #10 
a = 8'd131; b = 8'd57;  #10 
a = 8'd131; b = 8'd58;  #10 
a = 8'd131; b = 8'd59;  #10 
a = 8'd131; b = 8'd60;  #10 
a = 8'd131; b = 8'd61;  #10 
a = 8'd131; b = 8'd62;  #10 
a = 8'd131; b = 8'd63;  #10 
a = 8'd131; b = 8'd64;  #10 
a = 8'd131; b = 8'd65;  #10 
a = 8'd131; b = 8'd66;  #10 
a = 8'd131; b = 8'd67;  #10 
a = 8'd131; b = 8'd68;  #10 
a = 8'd131; b = 8'd69;  #10 
a = 8'd131; b = 8'd70;  #10 
a = 8'd131; b = 8'd71;  #10 
a = 8'd131; b = 8'd72;  #10 
a = 8'd131; b = 8'd73;  #10 
a = 8'd131; b = 8'd74;  #10 
a = 8'd131; b = 8'd75;  #10 
a = 8'd131; b = 8'd76;  #10 
a = 8'd131; b = 8'd77;  #10 
a = 8'd131; b = 8'd78;  #10 
a = 8'd131; b = 8'd79;  #10 
a = 8'd131; b = 8'd80;  #10 
a = 8'd131; b = 8'd81;  #10 
a = 8'd131; b = 8'd82;  #10 
a = 8'd131; b = 8'd83;  #10 
a = 8'd131; b = 8'd84;  #10 
a = 8'd131; b = 8'd85;  #10 
a = 8'd131; b = 8'd86;  #10 
a = 8'd131; b = 8'd87;  #10 
a = 8'd131; b = 8'd88;  #10 
a = 8'd131; b = 8'd89;  #10 
a = 8'd131; b = 8'd90;  #10 
a = 8'd131; b = 8'd91;  #10 
a = 8'd131; b = 8'd92;  #10 
a = 8'd131; b = 8'd93;  #10 
a = 8'd131; b = 8'd94;  #10 
a = 8'd131; b = 8'd95;  #10 
a = 8'd131; b = 8'd96;  #10 
a = 8'd131; b = 8'd97;  #10 
a = 8'd131; b = 8'd98;  #10 
a = 8'd131; b = 8'd99;  #10 
a = 8'd131; b = 8'd100;  #10 
a = 8'd131; b = 8'd101;  #10 
a = 8'd131; b = 8'd102;  #10 
a = 8'd131; b = 8'd103;  #10 
a = 8'd131; b = 8'd104;  #10 
a = 8'd131; b = 8'd105;  #10 
a = 8'd131; b = 8'd106;  #10 
a = 8'd131; b = 8'd107;  #10 
a = 8'd131; b = 8'd108;  #10 
a = 8'd131; b = 8'd109;  #10 
a = 8'd131; b = 8'd110;  #10 
a = 8'd131; b = 8'd111;  #10 
a = 8'd131; b = 8'd112;  #10 
a = 8'd131; b = 8'd113;  #10 
a = 8'd131; b = 8'd114;  #10 
a = 8'd131; b = 8'd115;  #10 
a = 8'd131; b = 8'd116;  #10 
a = 8'd131; b = 8'd117;  #10 
a = 8'd131; b = 8'd118;  #10 
a = 8'd131; b = 8'd119;  #10 
a = 8'd131; b = 8'd120;  #10 
a = 8'd131; b = 8'd121;  #10 
a = 8'd131; b = 8'd122;  #10 
a = 8'd131; b = 8'd123;  #10 
a = 8'd131; b = 8'd124;  #10 
a = 8'd131; b = 8'd125;  #10 
a = 8'd131; b = 8'd126;  #10 
a = 8'd131; b = 8'd127;  #10 
a = 8'd131; b = 8'd128;  #10 
a = 8'd131; b = 8'd129;  #10 
a = 8'd131; b = 8'd130;  #10 
a = 8'd131; b = 8'd131;  #10 
a = 8'd131; b = 8'd132;  #10 
a = 8'd131; b = 8'd133;  #10 
a = 8'd131; b = 8'd134;  #10 
a = 8'd131; b = 8'd135;  #10 
a = 8'd131; b = 8'd136;  #10 
a = 8'd131; b = 8'd137;  #10 
a = 8'd131; b = 8'd138;  #10 
a = 8'd131; b = 8'd139;  #10 
a = 8'd131; b = 8'd140;  #10 
a = 8'd131; b = 8'd141;  #10 
a = 8'd131; b = 8'd142;  #10 
a = 8'd131; b = 8'd143;  #10 
a = 8'd131; b = 8'd144;  #10 
a = 8'd131; b = 8'd145;  #10 
a = 8'd131; b = 8'd146;  #10 
a = 8'd131; b = 8'd147;  #10 
a = 8'd131; b = 8'd148;  #10 
a = 8'd131; b = 8'd149;  #10 
a = 8'd131; b = 8'd150;  #10 
a = 8'd131; b = 8'd151;  #10 
a = 8'd131; b = 8'd152;  #10 
a = 8'd131; b = 8'd153;  #10 
a = 8'd131; b = 8'd154;  #10 
a = 8'd131; b = 8'd155;  #10 
a = 8'd131; b = 8'd156;  #10 
a = 8'd131; b = 8'd157;  #10 
a = 8'd131; b = 8'd158;  #10 
a = 8'd131; b = 8'd159;  #10 
a = 8'd131; b = 8'd160;  #10 
a = 8'd131; b = 8'd161;  #10 
a = 8'd131; b = 8'd162;  #10 
a = 8'd131; b = 8'd163;  #10 
a = 8'd131; b = 8'd164;  #10 
a = 8'd131; b = 8'd165;  #10 
a = 8'd131; b = 8'd166;  #10 
a = 8'd131; b = 8'd167;  #10 
a = 8'd131; b = 8'd168;  #10 
a = 8'd131; b = 8'd169;  #10 
a = 8'd131; b = 8'd170;  #10 
a = 8'd131; b = 8'd171;  #10 
a = 8'd131; b = 8'd172;  #10 
a = 8'd131; b = 8'd173;  #10 
a = 8'd131; b = 8'd174;  #10 
a = 8'd131; b = 8'd175;  #10 
a = 8'd131; b = 8'd176;  #10 
a = 8'd131; b = 8'd177;  #10 
a = 8'd131; b = 8'd178;  #10 
a = 8'd131; b = 8'd179;  #10 
a = 8'd131; b = 8'd180;  #10 
a = 8'd131; b = 8'd181;  #10 
a = 8'd131; b = 8'd182;  #10 
a = 8'd131; b = 8'd183;  #10 
a = 8'd131; b = 8'd184;  #10 
a = 8'd131; b = 8'd185;  #10 
a = 8'd131; b = 8'd186;  #10 
a = 8'd131; b = 8'd187;  #10 
a = 8'd131; b = 8'd188;  #10 
a = 8'd131; b = 8'd189;  #10 
a = 8'd131; b = 8'd190;  #10 
a = 8'd131; b = 8'd191;  #10 
a = 8'd131; b = 8'd192;  #10 
a = 8'd131; b = 8'd193;  #10 
a = 8'd131; b = 8'd194;  #10 
a = 8'd131; b = 8'd195;  #10 
a = 8'd131; b = 8'd196;  #10 
a = 8'd131; b = 8'd197;  #10 
a = 8'd131; b = 8'd198;  #10 
a = 8'd131; b = 8'd199;  #10 
a = 8'd131; b = 8'd200;  #10 
a = 8'd131; b = 8'd201;  #10 
a = 8'd131; b = 8'd202;  #10 
a = 8'd131; b = 8'd203;  #10 
a = 8'd131; b = 8'd204;  #10 
a = 8'd131; b = 8'd205;  #10 
a = 8'd131; b = 8'd206;  #10 
a = 8'd131; b = 8'd207;  #10 
a = 8'd131; b = 8'd208;  #10 
a = 8'd131; b = 8'd209;  #10 
a = 8'd131; b = 8'd210;  #10 
a = 8'd131; b = 8'd211;  #10 
a = 8'd131; b = 8'd212;  #10 
a = 8'd131; b = 8'd213;  #10 
a = 8'd131; b = 8'd214;  #10 
a = 8'd131; b = 8'd215;  #10 
a = 8'd131; b = 8'd216;  #10 
a = 8'd131; b = 8'd217;  #10 
a = 8'd131; b = 8'd218;  #10 
a = 8'd131; b = 8'd219;  #10 
a = 8'd131; b = 8'd220;  #10 
a = 8'd131; b = 8'd221;  #10 
a = 8'd131; b = 8'd222;  #10 
a = 8'd131; b = 8'd223;  #10 
a = 8'd131; b = 8'd224;  #10 
a = 8'd131; b = 8'd225;  #10 
a = 8'd131; b = 8'd226;  #10 
a = 8'd131; b = 8'd227;  #10 
a = 8'd131; b = 8'd228;  #10 
a = 8'd131; b = 8'd229;  #10 
a = 8'd131; b = 8'd230;  #10 
a = 8'd131; b = 8'd231;  #10 
a = 8'd131; b = 8'd232;  #10 
a = 8'd131; b = 8'd233;  #10 
a = 8'd131; b = 8'd234;  #10 
a = 8'd131; b = 8'd235;  #10 
a = 8'd131; b = 8'd236;  #10 
a = 8'd131; b = 8'd237;  #10 
a = 8'd131; b = 8'd238;  #10 
a = 8'd131; b = 8'd239;  #10 
a = 8'd131; b = 8'd240;  #10 
a = 8'd131; b = 8'd241;  #10 
a = 8'd131; b = 8'd242;  #10 
a = 8'd131; b = 8'd243;  #10 
a = 8'd131; b = 8'd244;  #10 
a = 8'd131; b = 8'd245;  #10 
a = 8'd131; b = 8'd246;  #10 
a = 8'd131; b = 8'd247;  #10 
a = 8'd131; b = 8'd248;  #10 
a = 8'd131; b = 8'd249;  #10 
a = 8'd131; b = 8'd250;  #10 
a = 8'd131; b = 8'd251;  #10 
a = 8'd131; b = 8'd252;  #10 
a = 8'd131; b = 8'd253;  #10 
a = 8'd131; b = 8'd254;  #10 
a = 8'd131; b = 8'd255;  #10 
a = 8'd132; b = 8'd0;  #10 
a = 8'd132; b = 8'd1;  #10 
a = 8'd132; b = 8'd2;  #10 
a = 8'd132; b = 8'd3;  #10 
a = 8'd132; b = 8'd4;  #10 
a = 8'd132; b = 8'd5;  #10 
a = 8'd132; b = 8'd6;  #10 
a = 8'd132; b = 8'd7;  #10 
a = 8'd132; b = 8'd8;  #10 
a = 8'd132; b = 8'd9;  #10 
a = 8'd132; b = 8'd10;  #10 
a = 8'd132; b = 8'd11;  #10 
a = 8'd132; b = 8'd12;  #10 
a = 8'd132; b = 8'd13;  #10 
a = 8'd132; b = 8'd14;  #10 
a = 8'd132; b = 8'd15;  #10 
a = 8'd132; b = 8'd16;  #10 
a = 8'd132; b = 8'd17;  #10 
a = 8'd132; b = 8'd18;  #10 
a = 8'd132; b = 8'd19;  #10 
a = 8'd132; b = 8'd20;  #10 
a = 8'd132; b = 8'd21;  #10 
a = 8'd132; b = 8'd22;  #10 
a = 8'd132; b = 8'd23;  #10 
a = 8'd132; b = 8'd24;  #10 
a = 8'd132; b = 8'd25;  #10 
a = 8'd132; b = 8'd26;  #10 
a = 8'd132; b = 8'd27;  #10 
a = 8'd132; b = 8'd28;  #10 
a = 8'd132; b = 8'd29;  #10 
a = 8'd132; b = 8'd30;  #10 
a = 8'd132; b = 8'd31;  #10 
a = 8'd132; b = 8'd32;  #10 
a = 8'd132; b = 8'd33;  #10 
a = 8'd132; b = 8'd34;  #10 
a = 8'd132; b = 8'd35;  #10 
a = 8'd132; b = 8'd36;  #10 
a = 8'd132; b = 8'd37;  #10 
a = 8'd132; b = 8'd38;  #10 
a = 8'd132; b = 8'd39;  #10 
a = 8'd132; b = 8'd40;  #10 
a = 8'd132; b = 8'd41;  #10 
a = 8'd132; b = 8'd42;  #10 
a = 8'd132; b = 8'd43;  #10 
a = 8'd132; b = 8'd44;  #10 
a = 8'd132; b = 8'd45;  #10 
a = 8'd132; b = 8'd46;  #10 
a = 8'd132; b = 8'd47;  #10 
a = 8'd132; b = 8'd48;  #10 
a = 8'd132; b = 8'd49;  #10 
a = 8'd132; b = 8'd50;  #10 
a = 8'd132; b = 8'd51;  #10 
a = 8'd132; b = 8'd52;  #10 
a = 8'd132; b = 8'd53;  #10 
a = 8'd132; b = 8'd54;  #10 
a = 8'd132; b = 8'd55;  #10 
a = 8'd132; b = 8'd56;  #10 
a = 8'd132; b = 8'd57;  #10 
a = 8'd132; b = 8'd58;  #10 
a = 8'd132; b = 8'd59;  #10 
a = 8'd132; b = 8'd60;  #10 
a = 8'd132; b = 8'd61;  #10 
a = 8'd132; b = 8'd62;  #10 
a = 8'd132; b = 8'd63;  #10 
a = 8'd132; b = 8'd64;  #10 
a = 8'd132; b = 8'd65;  #10 
a = 8'd132; b = 8'd66;  #10 
a = 8'd132; b = 8'd67;  #10 
a = 8'd132; b = 8'd68;  #10 
a = 8'd132; b = 8'd69;  #10 
a = 8'd132; b = 8'd70;  #10 
a = 8'd132; b = 8'd71;  #10 
a = 8'd132; b = 8'd72;  #10 
a = 8'd132; b = 8'd73;  #10 
a = 8'd132; b = 8'd74;  #10 
a = 8'd132; b = 8'd75;  #10 
a = 8'd132; b = 8'd76;  #10 
a = 8'd132; b = 8'd77;  #10 
a = 8'd132; b = 8'd78;  #10 
a = 8'd132; b = 8'd79;  #10 
a = 8'd132; b = 8'd80;  #10 
a = 8'd132; b = 8'd81;  #10 
a = 8'd132; b = 8'd82;  #10 
a = 8'd132; b = 8'd83;  #10 
a = 8'd132; b = 8'd84;  #10 
a = 8'd132; b = 8'd85;  #10 
a = 8'd132; b = 8'd86;  #10 
a = 8'd132; b = 8'd87;  #10 
a = 8'd132; b = 8'd88;  #10 
a = 8'd132; b = 8'd89;  #10 
a = 8'd132; b = 8'd90;  #10 
a = 8'd132; b = 8'd91;  #10 
a = 8'd132; b = 8'd92;  #10 
a = 8'd132; b = 8'd93;  #10 
a = 8'd132; b = 8'd94;  #10 
a = 8'd132; b = 8'd95;  #10 
a = 8'd132; b = 8'd96;  #10 
a = 8'd132; b = 8'd97;  #10 
a = 8'd132; b = 8'd98;  #10 
a = 8'd132; b = 8'd99;  #10 
a = 8'd132; b = 8'd100;  #10 
a = 8'd132; b = 8'd101;  #10 
a = 8'd132; b = 8'd102;  #10 
a = 8'd132; b = 8'd103;  #10 
a = 8'd132; b = 8'd104;  #10 
a = 8'd132; b = 8'd105;  #10 
a = 8'd132; b = 8'd106;  #10 
a = 8'd132; b = 8'd107;  #10 
a = 8'd132; b = 8'd108;  #10 
a = 8'd132; b = 8'd109;  #10 
a = 8'd132; b = 8'd110;  #10 
a = 8'd132; b = 8'd111;  #10 
a = 8'd132; b = 8'd112;  #10 
a = 8'd132; b = 8'd113;  #10 
a = 8'd132; b = 8'd114;  #10 
a = 8'd132; b = 8'd115;  #10 
a = 8'd132; b = 8'd116;  #10 
a = 8'd132; b = 8'd117;  #10 
a = 8'd132; b = 8'd118;  #10 
a = 8'd132; b = 8'd119;  #10 
a = 8'd132; b = 8'd120;  #10 
a = 8'd132; b = 8'd121;  #10 
a = 8'd132; b = 8'd122;  #10 
a = 8'd132; b = 8'd123;  #10 
a = 8'd132; b = 8'd124;  #10 
a = 8'd132; b = 8'd125;  #10 
a = 8'd132; b = 8'd126;  #10 
a = 8'd132; b = 8'd127;  #10 
a = 8'd132; b = 8'd128;  #10 
a = 8'd132; b = 8'd129;  #10 
a = 8'd132; b = 8'd130;  #10 
a = 8'd132; b = 8'd131;  #10 
a = 8'd132; b = 8'd132;  #10 
a = 8'd132; b = 8'd133;  #10 
a = 8'd132; b = 8'd134;  #10 
a = 8'd132; b = 8'd135;  #10 
a = 8'd132; b = 8'd136;  #10 
a = 8'd132; b = 8'd137;  #10 
a = 8'd132; b = 8'd138;  #10 
a = 8'd132; b = 8'd139;  #10 
a = 8'd132; b = 8'd140;  #10 
a = 8'd132; b = 8'd141;  #10 
a = 8'd132; b = 8'd142;  #10 
a = 8'd132; b = 8'd143;  #10 
a = 8'd132; b = 8'd144;  #10 
a = 8'd132; b = 8'd145;  #10 
a = 8'd132; b = 8'd146;  #10 
a = 8'd132; b = 8'd147;  #10 
a = 8'd132; b = 8'd148;  #10 
a = 8'd132; b = 8'd149;  #10 
a = 8'd132; b = 8'd150;  #10 
a = 8'd132; b = 8'd151;  #10 
a = 8'd132; b = 8'd152;  #10 
a = 8'd132; b = 8'd153;  #10 
a = 8'd132; b = 8'd154;  #10 
a = 8'd132; b = 8'd155;  #10 
a = 8'd132; b = 8'd156;  #10 
a = 8'd132; b = 8'd157;  #10 
a = 8'd132; b = 8'd158;  #10 
a = 8'd132; b = 8'd159;  #10 
a = 8'd132; b = 8'd160;  #10 
a = 8'd132; b = 8'd161;  #10 
a = 8'd132; b = 8'd162;  #10 
a = 8'd132; b = 8'd163;  #10 
a = 8'd132; b = 8'd164;  #10 
a = 8'd132; b = 8'd165;  #10 
a = 8'd132; b = 8'd166;  #10 
a = 8'd132; b = 8'd167;  #10 
a = 8'd132; b = 8'd168;  #10 
a = 8'd132; b = 8'd169;  #10 
a = 8'd132; b = 8'd170;  #10 
a = 8'd132; b = 8'd171;  #10 
a = 8'd132; b = 8'd172;  #10 
a = 8'd132; b = 8'd173;  #10 
a = 8'd132; b = 8'd174;  #10 
a = 8'd132; b = 8'd175;  #10 
a = 8'd132; b = 8'd176;  #10 
a = 8'd132; b = 8'd177;  #10 
a = 8'd132; b = 8'd178;  #10 
a = 8'd132; b = 8'd179;  #10 
a = 8'd132; b = 8'd180;  #10 
a = 8'd132; b = 8'd181;  #10 
a = 8'd132; b = 8'd182;  #10 
a = 8'd132; b = 8'd183;  #10 
a = 8'd132; b = 8'd184;  #10 
a = 8'd132; b = 8'd185;  #10 
a = 8'd132; b = 8'd186;  #10 
a = 8'd132; b = 8'd187;  #10 
a = 8'd132; b = 8'd188;  #10 
a = 8'd132; b = 8'd189;  #10 
a = 8'd132; b = 8'd190;  #10 
a = 8'd132; b = 8'd191;  #10 
a = 8'd132; b = 8'd192;  #10 
a = 8'd132; b = 8'd193;  #10 
a = 8'd132; b = 8'd194;  #10 
a = 8'd132; b = 8'd195;  #10 
a = 8'd132; b = 8'd196;  #10 
a = 8'd132; b = 8'd197;  #10 
a = 8'd132; b = 8'd198;  #10 
a = 8'd132; b = 8'd199;  #10 
a = 8'd132; b = 8'd200;  #10 
a = 8'd132; b = 8'd201;  #10 
a = 8'd132; b = 8'd202;  #10 
a = 8'd132; b = 8'd203;  #10 
a = 8'd132; b = 8'd204;  #10 
a = 8'd132; b = 8'd205;  #10 
a = 8'd132; b = 8'd206;  #10 
a = 8'd132; b = 8'd207;  #10 
a = 8'd132; b = 8'd208;  #10 
a = 8'd132; b = 8'd209;  #10 
a = 8'd132; b = 8'd210;  #10 
a = 8'd132; b = 8'd211;  #10 
a = 8'd132; b = 8'd212;  #10 
a = 8'd132; b = 8'd213;  #10 
a = 8'd132; b = 8'd214;  #10 
a = 8'd132; b = 8'd215;  #10 
a = 8'd132; b = 8'd216;  #10 
a = 8'd132; b = 8'd217;  #10 
a = 8'd132; b = 8'd218;  #10 
a = 8'd132; b = 8'd219;  #10 
a = 8'd132; b = 8'd220;  #10 
a = 8'd132; b = 8'd221;  #10 
a = 8'd132; b = 8'd222;  #10 
a = 8'd132; b = 8'd223;  #10 
a = 8'd132; b = 8'd224;  #10 
a = 8'd132; b = 8'd225;  #10 
a = 8'd132; b = 8'd226;  #10 
a = 8'd132; b = 8'd227;  #10 
a = 8'd132; b = 8'd228;  #10 
a = 8'd132; b = 8'd229;  #10 
a = 8'd132; b = 8'd230;  #10 
a = 8'd132; b = 8'd231;  #10 
a = 8'd132; b = 8'd232;  #10 
a = 8'd132; b = 8'd233;  #10 
a = 8'd132; b = 8'd234;  #10 
a = 8'd132; b = 8'd235;  #10 
a = 8'd132; b = 8'd236;  #10 
a = 8'd132; b = 8'd237;  #10 
a = 8'd132; b = 8'd238;  #10 
a = 8'd132; b = 8'd239;  #10 
a = 8'd132; b = 8'd240;  #10 
a = 8'd132; b = 8'd241;  #10 
a = 8'd132; b = 8'd242;  #10 
a = 8'd132; b = 8'd243;  #10 
a = 8'd132; b = 8'd244;  #10 
a = 8'd132; b = 8'd245;  #10 
a = 8'd132; b = 8'd246;  #10 
a = 8'd132; b = 8'd247;  #10 
a = 8'd132; b = 8'd248;  #10 
a = 8'd132; b = 8'd249;  #10 
a = 8'd132; b = 8'd250;  #10 
a = 8'd132; b = 8'd251;  #10 
a = 8'd132; b = 8'd252;  #10 
a = 8'd132; b = 8'd253;  #10 
a = 8'd132; b = 8'd254;  #10 
a = 8'd132; b = 8'd255;  #10 
a = 8'd133; b = 8'd0;  #10 
a = 8'd133; b = 8'd1;  #10 
a = 8'd133; b = 8'd2;  #10 
a = 8'd133; b = 8'd3;  #10 
a = 8'd133; b = 8'd4;  #10 
a = 8'd133; b = 8'd5;  #10 
a = 8'd133; b = 8'd6;  #10 
a = 8'd133; b = 8'd7;  #10 
a = 8'd133; b = 8'd8;  #10 
a = 8'd133; b = 8'd9;  #10 
a = 8'd133; b = 8'd10;  #10 
a = 8'd133; b = 8'd11;  #10 
a = 8'd133; b = 8'd12;  #10 
a = 8'd133; b = 8'd13;  #10 
a = 8'd133; b = 8'd14;  #10 
a = 8'd133; b = 8'd15;  #10 
a = 8'd133; b = 8'd16;  #10 
a = 8'd133; b = 8'd17;  #10 
a = 8'd133; b = 8'd18;  #10 
a = 8'd133; b = 8'd19;  #10 
a = 8'd133; b = 8'd20;  #10 
a = 8'd133; b = 8'd21;  #10 
a = 8'd133; b = 8'd22;  #10 
a = 8'd133; b = 8'd23;  #10 
a = 8'd133; b = 8'd24;  #10 
a = 8'd133; b = 8'd25;  #10 
a = 8'd133; b = 8'd26;  #10 
a = 8'd133; b = 8'd27;  #10 
a = 8'd133; b = 8'd28;  #10 
a = 8'd133; b = 8'd29;  #10 
a = 8'd133; b = 8'd30;  #10 
a = 8'd133; b = 8'd31;  #10 
a = 8'd133; b = 8'd32;  #10 
a = 8'd133; b = 8'd33;  #10 
a = 8'd133; b = 8'd34;  #10 
a = 8'd133; b = 8'd35;  #10 
a = 8'd133; b = 8'd36;  #10 
a = 8'd133; b = 8'd37;  #10 
a = 8'd133; b = 8'd38;  #10 
a = 8'd133; b = 8'd39;  #10 
a = 8'd133; b = 8'd40;  #10 
a = 8'd133; b = 8'd41;  #10 
a = 8'd133; b = 8'd42;  #10 
a = 8'd133; b = 8'd43;  #10 
a = 8'd133; b = 8'd44;  #10 
a = 8'd133; b = 8'd45;  #10 
a = 8'd133; b = 8'd46;  #10 
a = 8'd133; b = 8'd47;  #10 
a = 8'd133; b = 8'd48;  #10 
a = 8'd133; b = 8'd49;  #10 
a = 8'd133; b = 8'd50;  #10 
a = 8'd133; b = 8'd51;  #10 
a = 8'd133; b = 8'd52;  #10 
a = 8'd133; b = 8'd53;  #10 
a = 8'd133; b = 8'd54;  #10 
a = 8'd133; b = 8'd55;  #10 
a = 8'd133; b = 8'd56;  #10 
a = 8'd133; b = 8'd57;  #10 
a = 8'd133; b = 8'd58;  #10 
a = 8'd133; b = 8'd59;  #10 
a = 8'd133; b = 8'd60;  #10 
a = 8'd133; b = 8'd61;  #10 
a = 8'd133; b = 8'd62;  #10 
a = 8'd133; b = 8'd63;  #10 
a = 8'd133; b = 8'd64;  #10 
a = 8'd133; b = 8'd65;  #10 
a = 8'd133; b = 8'd66;  #10 
a = 8'd133; b = 8'd67;  #10 
a = 8'd133; b = 8'd68;  #10 
a = 8'd133; b = 8'd69;  #10 
a = 8'd133; b = 8'd70;  #10 
a = 8'd133; b = 8'd71;  #10 
a = 8'd133; b = 8'd72;  #10 
a = 8'd133; b = 8'd73;  #10 
a = 8'd133; b = 8'd74;  #10 
a = 8'd133; b = 8'd75;  #10 
a = 8'd133; b = 8'd76;  #10 
a = 8'd133; b = 8'd77;  #10 
a = 8'd133; b = 8'd78;  #10 
a = 8'd133; b = 8'd79;  #10 
a = 8'd133; b = 8'd80;  #10 
a = 8'd133; b = 8'd81;  #10 
a = 8'd133; b = 8'd82;  #10 
a = 8'd133; b = 8'd83;  #10 
a = 8'd133; b = 8'd84;  #10 
a = 8'd133; b = 8'd85;  #10 
a = 8'd133; b = 8'd86;  #10 
a = 8'd133; b = 8'd87;  #10 
a = 8'd133; b = 8'd88;  #10 
a = 8'd133; b = 8'd89;  #10 
a = 8'd133; b = 8'd90;  #10 
a = 8'd133; b = 8'd91;  #10 
a = 8'd133; b = 8'd92;  #10 
a = 8'd133; b = 8'd93;  #10 
a = 8'd133; b = 8'd94;  #10 
a = 8'd133; b = 8'd95;  #10 
a = 8'd133; b = 8'd96;  #10 
a = 8'd133; b = 8'd97;  #10 
a = 8'd133; b = 8'd98;  #10 
a = 8'd133; b = 8'd99;  #10 
a = 8'd133; b = 8'd100;  #10 
a = 8'd133; b = 8'd101;  #10 
a = 8'd133; b = 8'd102;  #10 
a = 8'd133; b = 8'd103;  #10 
a = 8'd133; b = 8'd104;  #10 
a = 8'd133; b = 8'd105;  #10 
a = 8'd133; b = 8'd106;  #10 
a = 8'd133; b = 8'd107;  #10 
a = 8'd133; b = 8'd108;  #10 
a = 8'd133; b = 8'd109;  #10 
a = 8'd133; b = 8'd110;  #10 
a = 8'd133; b = 8'd111;  #10 
a = 8'd133; b = 8'd112;  #10 
a = 8'd133; b = 8'd113;  #10 
a = 8'd133; b = 8'd114;  #10 
a = 8'd133; b = 8'd115;  #10 
a = 8'd133; b = 8'd116;  #10 
a = 8'd133; b = 8'd117;  #10 
a = 8'd133; b = 8'd118;  #10 
a = 8'd133; b = 8'd119;  #10 
a = 8'd133; b = 8'd120;  #10 
a = 8'd133; b = 8'd121;  #10 
a = 8'd133; b = 8'd122;  #10 
a = 8'd133; b = 8'd123;  #10 
a = 8'd133; b = 8'd124;  #10 
a = 8'd133; b = 8'd125;  #10 
a = 8'd133; b = 8'd126;  #10 
a = 8'd133; b = 8'd127;  #10 
a = 8'd133; b = 8'd128;  #10 
a = 8'd133; b = 8'd129;  #10 
a = 8'd133; b = 8'd130;  #10 
a = 8'd133; b = 8'd131;  #10 
a = 8'd133; b = 8'd132;  #10 
a = 8'd133; b = 8'd133;  #10 
a = 8'd133; b = 8'd134;  #10 
a = 8'd133; b = 8'd135;  #10 
a = 8'd133; b = 8'd136;  #10 
a = 8'd133; b = 8'd137;  #10 
a = 8'd133; b = 8'd138;  #10 
a = 8'd133; b = 8'd139;  #10 
a = 8'd133; b = 8'd140;  #10 
a = 8'd133; b = 8'd141;  #10 
a = 8'd133; b = 8'd142;  #10 
a = 8'd133; b = 8'd143;  #10 
a = 8'd133; b = 8'd144;  #10 
a = 8'd133; b = 8'd145;  #10 
a = 8'd133; b = 8'd146;  #10 
a = 8'd133; b = 8'd147;  #10 
a = 8'd133; b = 8'd148;  #10 
a = 8'd133; b = 8'd149;  #10 
a = 8'd133; b = 8'd150;  #10 
a = 8'd133; b = 8'd151;  #10 
a = 8'd133; b = 8'd152;  #10 
a = 8'd133; b = 8'd153;  #10 
a = 8'd133; b = 8'd154;  #10 
a = 8'd133; b = 8'd155;  #10 
a = 8'd133; b = 8'd156;  #10 
a = 8'd133; b = 8'd157;  #10 
a = 8'd133; b = 8'd158;  #10 
a = 8'd133; b = 8'd159;  #10 
a = 8'd133; b = 8'd160;  #10 
a = 8'd133; b = 8'd161;  #10 
a = 8'd133; b = 8'd162;  #10 
a = 8'd133; b = 8'd163;  #10 
a = 8'd133; b = 8'd164;  #10 
a = 8'd133; b = 8'd165;  #10 
a = 8'd133; b = 8'd166;  #10 
a = 8'd133; b = 8'd167;  #10 
a = 8'd133; b = 8'd168;  #10 
a = 8'd133; b = 8'd169;  #10 
a = 8'd133; b = 8'd170;  #10 
a = 8'd133; b = 8'd171;  #10 
a = 8'd133; b = 8'd172;  #10 
a = 8'd133; b = 8'd173;  #10 
a = 8'd133; b = 8'd174;  #10 
a = 8'd133; b = 8'd175;  #10 
a = 8'd133; b = 8'd176;  #10 
a = 8'd133; b = 8'd177;  #10 
a = 8'd133; b = 8'd178;  #10 
a = 8'd133; b = 8'd179;  #10 
a = 8'd133; b = 8'd180;  #10 
a = 8'd133; b = 8'd181;  #10 
a = 8'd133; b = 8'd182;  #10 
a = 8'd133; b = 8'd183;  #10 
a = 8'd133; b = 8'd184;  #10 
a = 8'd133; b = 8'd185;  #10 
a = 8'd133; b = 8'd186;  #10 
a = 8'd133; b = 8'd187;  #10 
a = 8'd133; b = 8'd188;  #10 
a = 8'd133; b = 8'd189;  #10 
a = 8'd133; b = 8'd190;  #10 
a = 8'd133; b = 8'd191;  #10 
a = 8'd133; b = 8'd192;  #10 
a = 8'd133; b = 8'd193;  #10 
a = 8'd133; b = 8'd194;  #10 
a = 8'd133; b = 8'd195;  #10 
a = 8'd133; b = 8'd196;  #10 
a = 8'd133; b = 8'd197;  #10 
a = 8'd133; b = 8'd198;  #10 
a = 8'd133; b = 8'd199;  #10 
a = 8'd133; b = 8'd200;  #10 
a = 8'd133; b = 8'd201;  #10 
a = 8'd133; b = 8'd202;  #10 
a = 8'd133; b = 8'd203;  #10 
a = 8'd133; b = 8'd204;  #10 
a = 8'd133; b = 8'd205;  #10 
a = 8'd133; b = 8'd206;  #10 
a = 8'd133; b = 8'd207;  #10 
a = 8'd133; b = 8'd208;  #10 
a = 8'd133; b = 8'd209;  #10 
a = 8'd133; b = 8'd210;  #10 
a = 8'd133; b = 8'd211;  #10 
a = 8'd133; b = 8'd212;  #10 
a = 8'd133; b = 8'd213;  #10 
a = 8'd133; b = 8'd214;  #10 
a = 8'd133; b = 8'd215;  #10 
a = 8'd133; b = 8'd216;  #10 
a = 8'd133; b = 8'd217;  #10 
a = 8'd133; b = 8'd218;  #10 
a = 8'd133; b = 8'd219;  #10 
a = 8'd133; b = 8'd220;  #10 
a = 8'd133; b = 8'd221;  #10 
a = 8'd133; b = 8'd222;  #10 
a = 8'd133; b = 8'd223;  #10 
a = 8'd133; b = 8'd224;  #10 
a = 8'd133; b = 8'd225;  #10 
a = 8'd133; b = 8'd226;  #10 
a = 8'd133; b = 8'd227;  #10 
a = 8'd133; b = 8'd228;  #10 
a = 8'd133; b = 8'd229;  #10 
a = 8'd133; b = 8'd230;  #10 
a = 8'd133; b = 8'd231;  #10 
a = 8'd133; b = 8'd232;  #10 
a = 8'd133; b = 8'd233;  #10 
a = 8'd133; b = 8'd234;  #10 
a = 8'd133; b = 8'd235;  #10 
a = 8'd133; b = 8'd236;  #10 
a = 8'd133; b = 8'd237;  #10 
a = 8'd133; b = 8'd238;  #10 
a = 8'd133; b = 8'd239;  #10 
a = 8'd133; b = 8'd240;  #10 
a = 8'd133; b = 8'd241;  #10 
a = 8'd133; b = 8'd242;  #10 
a = 8'd133; b = 8'd243;  #10 
a = 8'd133; b = 8'd244;  #10 
a = 8'd133; b = 8'd245;  #10 
a = 8'd133; b = 8'd246;  #10 
a = 8'd133; b = 8'd247;  #10 
a = 8'd133; b = 8'd248;  #10 
a = 8'd133; b = 8'd249;  #10 
a = 8'd133; b = 8'd250;  #10 
a = 8'd133; b = 8'd251;  #10 
a = 8'd133; b = 8'd252;  #10 
a = 8'd133; b = 8'd253;  #10 
a = 8'd133; b = 8'd254;  #10 
a = 8'd133; b = 8'd255;  #10 
a = 8'd134; b = 8'd0;  #10 
a = 8'd134; b = 8'd1;  #10 
a = 8'd134; b = 8'd2;  #10 
a = 8'd134; b = 8'd3;  #10 
a = 8'd134; b = 8'd4;  #10 
a = 8'd134; b = 8'd5;  #10 
a = 8'd134; b = 8'd6;  #10 
a = 8'd134; b = 8'd7;  #10 
a = 8'd134; b = 8'd8;  #10 
a = 8'd134; b = 8'd9;  #10 
a = 8'd134; b = 8'd10;  #10 
a = 8'd134; b = 8'd11;  #10 
a = 8'd134; b = 8'd12;  #10 
a = 8'd134; b = 8'd13;  #10 
a = 8'd134; b = 8'd14;  #10 
a = 8'd134; b = 8'd15;  #10 
a = 8'd134; b = 8'd16;  #10 
a = 8'd134; b = 8'd17;  #10 
a = 8'd134; b = 8'd18;  #10 
a = 8'd134; b = 8'd19;  #10 
a = 8'd134; b = 8'd20;  #10 
a = 8'd134; b = 8'd21;  #10 
a = 8'd134; b = 8'd22;  #10 
a = 8'd134; b = 8'd23;  #10 
a = 8'd134; b = 8'd24;  #10 
a = 8'd134; b = 8'd25;  #10 
a = 8'd134; b = 8'd26;  #10 
a = 8'd134; b = 8'd27;  #10 
a = 8'd134; b = 8'd28;  #10 
a = 8'd134; b = 8'd29;  #10 
a = 8'd134; b = 8'd30;  #10 
a = 8'd134; b = 8'd31;  #10 
a = 8'd134; b = 8'd32;  #10 
a = 8'd134; b = 8'd33;  #10 
a = 8'd134; b = 8'd34;  #10 
a = 8'd134; b = 8'd35;  #10 
a = 8'd134; b = 8'd36;  #10 
a = 8'd134; b = 8'd37;  #10 
a = 8'd134; b = 8'd38;  #10 
a = 8'd134; b = 8'd39;  #10 
a = 8'd134; b = 8'd40;  #10 
a = 8'd134; b = 8'd41;  #10 
a = 8'd134; b = 8'd42;  #10 
a = 8'd134; b = 8'd43;  #10 
a = 8'd134; b = 8'd44;  #10 
a = 8'd134; b = 8'd45;  #10 
a = 8'd134; b = 8'd46;  #10 
a = 8'd134; b = 8'd47;  #10 
a = 8'd134; b = 8'd48;  #10 
a = 8'd134; b = 8'd49;  #10 
a = 8'd134; b = 8'd50;  #10 
a = 8'd134; b = 8'd51;  #10 
a = 8'd134; b = 8'd52;  #10 
a = 8'd134; b = 8'd53;  #10 
a = 8'd134; b = 8'd54;  #10 
a = 8'd134; b = 8'd55;  #10 
a = 8'd134; b = 8'd56;  #10 
a = 8'd134; b = 8'd57;  #10 
a = 8'd134; b = 8'd58;  #10 
a = 8'd134; b = 8'd59;  #10 
a = 8'd134; b = 8'd60;  #10 
a = 8'd134; b = 8'd61;  #10 
a = 8'd134; b = 8'd62;  #10 
a = 8'd134; b = 8'd63;  #10 
a = 8'd134; b = 8'd64;  #10 
a = 8'd134; b = 8'd65;  #10 
a = 8'd134; b = 8'd66;  #10 
a = 8'd134; b = 8'd67;  #10 
a = 8'd134; b = 8'd68;  #10 
a = 8'd134; b = 8'd69;  #10 
a = 8'd134; b = 8'd70;  #10 
a = 8'd134; b = 8'd71;  #10 
a = 8'd134; b = 8'd72;  #10 
a = 8'd134; b = 8'd73;  #10 
a = 8'd134; b = 8'd74;  #10 
a = 8'd134; b = 8'd75;  #10 
a = 8'd134; b = 8'd76;  #10 
a = 8'd134; b = 8'd77;  #10 
a = 8'd134; b = 8'd78;  #10 
a = 8'd134; b = 8'd79;  #10 
a = 8'd134; b = 8'd80;  #10 
a = 8'd134; b = 8'd81;  #10 
a = 8'd134; b = 8'd82;  #10 
a = 8'd134; b = 8'd83;  #10 
a = 8'd134; b = 8'd84;  #10 
a = 8'd134; b = 8'd85;  #10 
a = 8'd134; b = 8'd86;  #10 
a = 8'd134; b = 8'd87;  #10 
a = 8'd134; b = 8'd88;  #10 
a = 8'd134; b = 8'd89;  #10 
a = 8'd134; b = 8'd90;  #10 
a = 8'd134; b = 8'd91;  #10 
a = 8'd134; b = 8'd92;  #10 
a = 8'd134; b = 8'd93;  #10 
a = 8'd134; b = 8'd94;  #10 
a = 8'd134; b = 8'd95;  #10 
a = 8'd134; b = 8'd96;  #10 
a = 8'd134; b = 8'd97;  #10 
a = 8'd134; b = 8'd98;  #10 
a = 8'd134; b = 8'd99;  #10 
a = 8'd134; b = 8'd100;  #10 
a = 8'd134; b = 8'd101;  #10 
a = 8'd134; b = 8'd102;  #10 
a = 8'd134; b = 8'd103;  #10 
a = 8'd134; b = 8'd104;  #10 
a = 8'd134; b = 8'd105;  #10 
a = 8'd134; b = 8'd106;  #10 
a = 8'd134; b = 8'd107;  #10 
a = 8'd134; b = 8'd108;  #10 
a = 8'd134; b = 8'd109;  #10 
a = 8'd134; b = 8'd110;  #10 
a = 8'd134; b = 8'd111;  #10 
a = 8'd134; b = 8'd112;  #10 
a = 8'd134; b = 8'd113;  #10 
a = 8'd134; b = 8'd114;  #10 
a = 8'd134; b = 8'd115;  #10 
a = 8'd134; b = 8'd116;  #10 
a = 8'd134; b = 8'd117;  #10 
a = 8'd134; b = 8'd118;  #10 
a = 8'd134; b = 8'd119;  #10 
a = 8'd134; b = 8'd120;  #10 
a = 8'd134; b = 8'd121;  #10 
a = 8'd134; b = 8'd122;  #10 
a = 8'd134; b = 8'd123;  #10 
a = 8'd134; b = 8'd124;  #10 
a = 8'd134; b = 8'd125;  #10 
a = 8'd134; b = 8'd126;  #10 
a = 8'd134; b = 8'd127;  #10 
a = 8'd134; b = 8'd128;  #10 
a = 8'd134; b = 8'd129;  #10 
a = 8'd134; b = 8'd130;  #10 
a = 8'd134; b = 8'd131;  #10 
a = 8'd134; b = 8'd132;  #10 
a = 8'd134; b = 8'd133;  #10 
a = 8'd134; b = 8'd134;  #10 
a = 8'd134; b = 8'd135;  #10 
a = 8'd134; b = 8'd136;  #10 
a = 8'd134; b = 8'd137;  #10 
a = 8'd134; b = 8'd138;  #10 
a = 8'd134; b = 8'd139;  #10 
a = 8'd134; b = 8'd140;  #10 
a = 8'd134; b = 8'd141;  #10 
a = 8'd134; b = 8'd142;  #10 
a = 8'd134; b = 8'd143;  #10 
a = 8'd134; b = 8'd144;  #10 
a = 8'd134; b = 8'd145;  #10 
a = 8'd134; b = 8'd146;  #10 
a = 8'd134; b = 8'd147;  #10 
a = 8'd134; b = 8'd148;  #10 
a = 8'd134; b = 8'd149;  #10 
a = 8'd134; b = 8'd150;  #10 
a = 8'd134; b = 8'd151;  #10 
a = 8'd134; b = 8'd152;  #10 
a = 8'd134; b = 8'd153;  #10 
a = 8'd134; b = 8'd154;  #10 
a = 8'd134; b = 8'd155;  #10 
a = 8'd134; b = 8'd156;  #10 
a = 8'd134; b = 8'd157;  #10 
a = 8'd134; b = 8'd158;  #10 
a = 8'd134; b = 8'd159;  #10 
a = 8'd134; b = 8'd160;  #10 
a = 8'd134; b = 8'd161;  #10 
a = 8'd134; b = 8'd162;  #10 
a = 8'd134; b = 8'd163;  #10 
a = 8'd134; b = 8'd164;  #10 
a = 8'd134; b = 8'd165;  #10 
a = 8'd134; b = 8'd166;  #10 
a = 8'd134; b = 8'd167;  #10 
a = 8'd134; b = 8'd168;  #10 
a = 8'd134; b = 8'd169;  #10 
a = 8'd134; b = 8'd170;  #10 
a = 8'd134; b = 8'd171;  #10 
a = 8'd134; b = 8'd172;  #10 
a = 8'd134; b = 8'd173;  #10 
a = 8'd134; b = 8'd174;  #10 
a = 8'd134; b = 8'd175;  #10 
a = 8'd134; b = 8'd176;  #10 
a = 8'd134; b = 8'd177;  #10 
a = 8'd134; b = 8'd178;  #10 
a = 8'd134; b = 8'd179;  #10 
a = 8'd134; b = 8'd180;  #10 
a = 8'd134; b = 8'd181;  #10 
a = 8'd134; b = 8'd182;  #10 
a = 8'd134; b = 8'd183;  #10 
a = 8'd134; b = 8'd184;  #10 
a = 8'd134; b = 8'd185;  #10 
a = 8'd134; b = 8'd186;  #10 
a = 8'd134; b = 8'd187;  #10 
a = 8'd134; b = 8'd188;  #10 
a = 8'd134; b = 8'd189;  #10 
a = 8'd134; b = 8'd190;  #10 
a = 8'd134; b = 8'd191;  #10 
a = 8'd134; b = 8'd192;  #10 
a = 8'd134; b = 8'd193;  #10 
a = 8'd134; b = 8'd194;  #10 
a = 8'd134; b = 8'd195;  #10 
a = 8'd134; b = 8'd196;  #10 
a = 8'd134; b = 8'd197;  #10 
a = 8'd134; b = 8'd198;  #10 
a = 8'd134; b = 8'd199;  #10 
a = 8'd134; b = 8'd200;  #10 
a = 8'd134; b = 8'd201;  #10 
a = 8'd134; b = 8'd202;  #10 
a = 8'd134; b = 8'd203;  #10 
a = 8'd134; b = 8'd204;  #10 
a = 8'd134; b = 8'd205;  #10 
a = 8'd134; b = 8'd206;  #10 
a = 8'd134; b = 8'd207;  #10 
a = 8'd134; b = 8'd208;  #10 
a = 8'd134; b = 8'd209;  #10 
a = 8'd134; b = 8'd210;  #10 
a = 8'd134; b = 8'd211;  #10 
a = 8'd134; b = 8'd212;  #10 
a = 8'd134; b = 8'd213;  #10 
a = 8'd134; b = 8'd214;  #10 
a = 8'd134; b = 8'd215;  #10 
a = 8'd134; b = 8'd216;  #10 
a = 8'd134; b = 8'd217;  #10 
a = 8'd134; b = 8'd218;  #10 
a = 8'd134; b = 8'd219;  #10 
a = 8'd134; b = 8'd220;  #10 
a = 8'd134; b = 8'd221;  #10 
a = 8'd134; b = 8'd222;  #10 
a = 8'd134; b = 8'd223;  #10 
a = 8'd134; b = 8'd224;  #10 
a = 8'd134; b = 8'd225;  #10 
a = 8'd134; b = 8'd226;  #10 
a = 8'd134; b = 8'd227;  #10 
a = 8'd134; b = 8'd228;  #10 
a = 8'd134; b = 8'd229;  #10 
a = 8'd134; b = 8'd230;  #10 
a = 8'd134; b = 8'd231;  #10 
a = 8'd134; b = 8'd232;  #10 
a = 8'd134; b = 8'd233;  #10 
a = 8'd134; b = 8'd234;  #10 
a = 8'd134; b = 8'd235;  #10 
a = 8'd134; b = 8'd236;  #10 
a = 8'd134; b = 8'd237;  #10 
a = 8'd134; b = 8'd238;  #10 
a = 8'd134; b = 8'd239;  #10 
a = 8'd134; b = 8'd240;  #10 
a = 8'd134; b = 8'd241;  #10 
a = 8'd134; b = 8'd242;  #10 
a = 8'd134; b = 8'd243;  #10 
a = 8'd134; b = 8'd244;  #10 
a = 8'd134; b = 8'd245;  #10 
a = 8'd134; b = 8'd246;  #10 
a = 8'd134; b = 8'd247;  #10 
a = 8'd134; b = 8'd248;  #10 
a = 8'd134; b = 8'd249;  #10 
a = 8'd134; b = 8'd250;  #10 
a = 8'd134; b = 8'd251;  #10 
a = 8'd134; b = 8'd252;  #10 
a = 8'd134; b = 8'd253;  #10 
a = 8'd134; b = 8'd254;  #10 
a = 8'd134; b = 8'd255;  #10 
a = 8'd135; b = 8'd0;  #10 
a = 8'd135; b = 8'd1;  #10 
a = 8'd135; b = 8'd2;  #10 
a = 8'd135; b = 8'd3;  #10 
a = 8'd135; b = 8'd4;  #10 
a = 8'd135; b = 8'd5;  #10 
a = 8'd135; b = 8'd6;  #10 
a = 8'd135; b = 8'd7;  #10 
a = 8'd135; b = 8'd8;  #10 
a = 8'd135; b = 8'd9;  #10 
a = 8'd135; b = 8'd10;  #10 
a = 8'd135; b = 8'd11;  #10 
a = 8'd135; b = 8'd12;  #10 
a = 8'd135; b = 8'd13;  #10 
a = 8'd135; b = 8'd14;  #10 
a = 8'd135; b = 8'd15;  #10 
a = 8'd135; b = 8'd16;  #10 
a = 8'd135; b = 8'd17;  #10 
a = 8'd135; b = 8'd18;  #10 
a = 8'd135; b = 8'd19;  #10 
a = 8'd135; b = 8'd20;  #10 
a = 8'd135; b = 8'd21;  #10 
a = 8'd135; b = 8'd22;  #10 
a = 8'd135; b = 8'd23;  #10 
a = 8'd135; b = 8'd24;  #10 
a = 8'd135; b = 8'd25;  #10 
a = 8'd135; b = 8'd26;  #10 
a = 8'd135; b = 8'd27;  #10 
a = 8'd135; b = 8'd28;  #10 
a = 8'd135; b = 8'd29;  #10 
a = 8'd135; b = 8'd30;  #10 
a = 8'd135; b = 8'd31;  #10 
a = 8'd135; b = 8'd32;  #10 
a = 8'd135; b = 8'd33;  #10 
a = 8'd135; b = 8'd34;  #10 
a = 8'd135; b = 8'd35;  #10 
a = 8'd135; b = 8'd36;  #10 
a = 8'd135; b = 8'd37;  #10 
a = 8'd135; b = 8'd38;  #10 
a = 8'd135; b = 8'd39;  #10 
a = 8'd135; b = 8'd40;  #10 
a = 8'd135; b = 8'd41;  #10 
a = 8'd135; b = 8'd42;  #10 
a = 8'd135; b = 8'd43;  #10 
a = 8'd135; b = 8'd44;  #10 
a = 8'd135; b = 8'd45;  #10 
a = 8'd135; b = 8'd46;  #10 
a = 8'd135; b = 8'd47;  #10 
a = 8'd135; b = 8'd48;  #10 
a = 8'd135; b = 8'd49;  #10 
a = 8'd135; b = 8'd50;  #10 
a = 8'd135; b = 8'd51;  #10 
a = 8'd135; b = 8'd52;  #10 
a = 8'd135; b = 8'd53;  #10 
a = 8'd135; b = 8'd54;  #10 
a = 8'd135; b = 8'd55;  #10 
a = 8'd135; b = 8'd56;  #10 
a = 8'd135; b = 8'd57;  #10 
a = 8'd135; b = 8'd58;  #10 
a = 8'd135; b = 8'd59;  #10 
a = 8'd135; b = 8'd60;  #10 
a = 8'd135; b = 8'd61;  #10 
a = 8'd135; b = 8'd62;  #10 
a = 8'd135; b = 8'd63;  #10 
a = 8'd135; b = 8'd64;  #10 
a = 8'd135; b = 8'd65;  #10 
a = 8'd135; b = 8'd66;  #10 
a = 8'd135; b = 8'd67;  #10 
a = 8'd135; b = 8'd68;  #10 
a = 8'd135; b = 8'd69;  #10 
a = 8'd135; b = 8'd70;  #10 
a = 8'd135; b = 8'd71;  #10 
a = 8'd135; b = 8'd72;  #10 
a = 8'd135; b = 8'd73;  #10 
a = 8'd135; b = 8'd74;  #10 
a = 8'd135; b = 8'd75;  #10 
a = 8'd135; b = 8'd76;  #10 
a = 8'd135; b = 8'd77;  #10 
a = 8'd135; b = 8'd78;  #10 
a = 8'd135; b = 8'd79;  #10 
a = 8'd135; b = 8'd80;  #10 
a = 8'd135; b = 8'd81;  #10 
a = 8'd135; b = 8'd82;  #10 
a = 8'd135; b = 8'd83;  #10 
a = 8'd135; b = 8'd84;  #10 
a = 8'd135; b = 8'd85;  #10 
a = 8'd135; b = 8'd86;  #10 
a = 8'd135; b = 8'd87;  #10 
a = 8'd135; b = 8'd88;  #10 
a = 8'd135; b = 8'd89;  #10 
a = 8'd135; b = 8'd90;  #10 
a = 8'd135; b = 8'd91;  #10 
a = 8'd135; b = 8'd92;  #10 
a = 8'd135; b = 8'd93;  #10 
a = 8'd135; b = 8'd94;  #10 
a = 8'd135; b = 8'd95;  #10 
a = 8'd135; b = 8'd96;  #10 
a = 8'd135; b = 8'd97;  #10 
a = 8'd135; b = 8'd98;  #10 
a = 8'd135; b = 8'd99;  #10 
a = 8'd135; b = 8'd100;  #10 
a = 8'd135; b = 8'd101;  #10 
a = 8'd135; b = 8'd102;  #10 
a = 8'd135; b = 8'd103;  #10 
a = 8'd135; b = 8'd104;  #10 
a = 8'd135; b = 8'd105;  #10 
a = 8'd135; b = 8'd106;  #10 
a = 8'd135; b = 8'd107;  #10 
a = 8'd135; b = 8'd108;  #10 
a = 8'd135; b = 8'd109;  #10 
a = 8'd135; b = 8'd110;  #10 
a = 8'd135; b = 8'd111;  #10 
a = 8'd135; b = 8'd112;  #10 
a = 8'd135; b = 8'd113;  #10 
a = 8'd135; b = 8'd114;  #10 
a = 8'd135; b = 8'd115;  #10 
a = 8'd135; b = 8'd116;  #10 
a = 8'd135; b = 8'd117;  #10 
a = 8'd135; b = 8'd118;  #10 
a = 8'd135; b = 8'd119;  #10 
a = 8'd135; b = 8'd120;  #10 
a = 8'd135; b = 8'd121;  #10 
a = 8'd135; b = 8'd122;  #10 
a = 8'd135; b = 8'd123;  #10 
a = 8'd135; b = 8'd124;  #10 
a = 8'd135; b = 8'd125;  #10 
a = 8'd135; b = 8'd126;  #10 
a = 8'd135; b = 8'd127;  #10 
a = 8'd135; b = 8'd128;  #10 
a = 8'd135; b = 8'd129;  #10 
a = 8'd135; b = 8'd130;  #10 
a = 8'd135; b = 8'd131;  #10 
a = 8'd135; b = 8'd132;  #10 
a = 8'd135; b = 8'd133;  #10 
a = 8'd135; b = 8'd134;  #10 
a = 8'd135; b = 8'd135;  #10 
a = 8'd135; b = 8'd136;  #10 
a = 8'd135; b = 8'd137;  #10 
a = 8'd135; b = 8'd138;  #10 
a = 8'd135; b = 8'd139;  #10 
a = 8'd135; b = 8'd140;  #10 
a = 8'd135; b = 8'd141;  #10 
a = 8'd135; b = 8'd142;  #10 
a = 8'd135; b = 8'd143;  #10 
a = 8'd135; b = 8'd144;  #10 
a = 8'd135; b = 8'd145;  #10 
a = 8'd135; b = 8'd146;  #10 
a = 8'd135; b = 8'd147;  #10 
a = 8'd135; b = 8'd148;  #10 
a = 8'd135; b = 8'd149;  #10 
a = 8'd135; b = 8'd150;  #10 
a = 8'd135; b = 8'd151;  #10 
a = 8'd135; b = 8'd152;  #10 
a = 8'd135; b = 8'd153;  #10 
a = 8'd135; b = 8'd154;  #10 
a = 8'd135; b = 8'd155;  #10 
a = 8'd135; b = 8'd156;  #10 
a = 8'd135; b = 8'd157;  #10 
a = 8'd135; b = 8'd158;  #10 
a = 8'd135; b = 8'd159;  #10 
a = 8'd135; b = 8'd160;  #10 
a = 8'd135; b = 8'd161;  #10 
a = 8'd135; b = 8'd162;  #10 
a = 8'd135; b = 8'd163;  #10 
a = 8'd135; b = 8'd164;  #10 
a = 8'd135; b = 8'd165;  #10 
a = 8'd135; b = 8'd166;  #10 
a = 8'd135; b = 8'd167;  #10 
a = 8'd135; b = 8'd168;  #10 
a = 8'd135; b = 8'd169;  #10 
a = 8'd135; b = 8'd170;  #10 
a = 8'd135; b = 8'd171;  #10 
a = 8'd135; b = 8'd172;  #10 
a = 8'd135; b = 8'd173;  #10 
a = 8'd135; b = 8'd174;  #10 
a = 8'd135; b = 8'd175;  #10 
a = 8'd135; b = 8'd176;  #10 
a = 8'd135; b = 8'd177;  #10 
a = 8'd135; b = 8'd178;  #10 
a = 8'd135; b = 8'd179;  #10 
a = 8'd135; b = 8'd180;  #10 
a = 8'd135; b = 8'd181;  #10 
a = 8'd135; b = 8'd182;  #10 
a = 8'd135; b = 8'd183;  #10 
a = 8'd135; b = 8'd184;  #10 
a = 8'd135; b = 8'd185;  #10 
a = 8'd135; b = 8'd186;  #10 
a = 8'd135; b = 8'd187;  #10 
a = 8'd135; b = 8'd188;  #10 
a = 8'd135; b = 8'd189;  #10 
a = 8'd135; b = 8'd190;  #10 
a = 8'd135; b = 8'd191;  #10 
a = 8'd135; b = 8'd192;  #10 
a = 8'd135; b = 8'd193;  #10 
a = 8'd135; b = 8'd194;  #10 
a = 8'd135; b = 8'd195;  #10 
a = 8'd135; b = 8'd196;  #10 
a = 8'd135; b = 8'd197;  #10 
a = 8'd135; b = 8'd198;  #10 
a = 8'd135; b = 8'd199;  #10 
a = 8'd135; b = 8'd200;  #10 
a = 8'd135; b = 8'd201;  #10 
a = 8'd135; b = 8'd202;  #10 
a = 8'd135; b = 8'd203;  #10 
a = 8'd135; b = 8'd204;  #10 
a = 8'd135; b = 8'd205;  #10 
a = 8'd135; b = 8'd206;  #10 
a = 8'd135; b = 8'd207;  #10 
a = 8'd135; b = 8'd208;  #10 
a = 8'd135; b = 8'd209;  #10 
a = 8'd135; b = 8'd210;  #10 
a = 8'd135; b = 8'd211;  #10 
a = 8'd135; b = 8'd212;  #10 
a = 8'd135; b = 8'd213;  #10 
a = 8'd135; b = 8'd214;  #10 
a = 8'd135; b = 8'd215;  #10 
a = 8'd135; b = 8'd216;  #10 
a = 8'd135; b = 8'd217;  #10 
a = 8'd135; b = 8'd218;  #10 
a = 8'd135; b = 8'd219;  #10 
a = 8'd135; b = 8'd220;  #10 
a = 8'd135; b = 8'd221;  #10 
a = 8'd135; b = 8'd222;  #10 
a = 8'd135; b = 8'd223;  #10 
a = 8'd135; b = 8'd224;  #10 
a = 8'd135; b = 8'd225;  #10 
a = 8'd135; b = 8'd226;  #10 
a = 8'd135; b = 8'd227;  #10 
a = 8'd135; b = 8'd228;  #10 
a = 8'd135; b = 8'd229;  #10 
a = 8'd135; b = 8'd230;  #10 
a = 8'd135; b = 8'd231;  #10 
a = 8'd135; b = 8'd232;  #10 
a = 8'd135; b = 8'd233;  #10 
a = 8'd135; b = 8'd234;  #10 
a = 8'd135; b = 8'd235;  #10 
a = 8'd135; b = 8'd236;  #10 
a = 8'd135; b = 8'd237;  #10 
a = 8'd135; b = 8'd238;  #10 
a = 8'd135; b = 8'd239;  #10 
a = 8'd135; b = 8'd240;  #10 
a = 8'd135; b = 8'd241;  #10 
a = 8'd135; b = 8'd242;  #10 
a = 8'd135; b = 8'd243;  #10 
a = 8'd135; b = 8'd244;  #10 
a = 8'd135; b = 8'd245;  #10 
a = 8'd135; b = 8'd246;  #10 
a = 8'd135; b = 8'd247;  #10 
a = 8'd135; b = 8'd248;  #10 
a = 8'd135; b = 8'd249;  #10 
a = 8'd135; b = 8'd250;  #10 
a = 8'd135; b = 8'd251;  #10 
a = 8'd135; b = 8'd252;  #10 
a = 8'd135; b = 8'd253;  #10 
a = 8'd135; b = 8'd254;  #10 
a = 8'd135; b = 8'd255;  #10 
a = 8'd136; b = 8'd0;  #10 
a = 8'd136; b = 8'd1;  #10 
a = 8'd136; b = 8'd2;  #10 
a = 8'd136; b = 8'd3;  #10 
a = 8'd136; b = 8'd4;  #10 
a = 8'd136; b = 8'd5;  #10 
a = 8'd136; b = 8'd6;  #10 
a = 8'd136; b = 8'd7;  #10 
a = 8'd136; b = 8'd8;  #10 
a = 8'd136; b = 8'd9;  #10 
a = 8'd136; b = 8'd10;  #10 
a = 8'd136; b = 8'd11;  #10 
a = 8'd136; b = 8'd12;  #10 
a = 8'd136; b = 8'd13;  #10 
a = 8'd136; b = 8'd14;  #10 
a = 8'd136; b = 8'd15;  #10 
a = 8'd136; b = 8'd16;  #10 
a = 8'd136; b = 8'd17;  #10 
a = 8'd136; b = 8'd18;  #10 
a = 8'd136; b = 8'd19;  #10 
a = 8'd136; b = 8'd20;  #10 
a = 8'd136; b = 8'd21;  #10 
a = 8'd136; b = 8'd22;  #10 
a = 8'd136; b = 8'd23;  #10 
a = 8'd136; b = 8'd24;  #10 
a = 8'd136; b = 8'd25;  #10 
a = 8'd136; b = 8'd26;  #10 
a = 8'd136; b = 8'd27;  #10 
a = 8'd136; b = 8'd28;  #10 
a = 8'd136; b = 8'd29;  #10 
a = 8'd136; b = 8'd30;  #10 
a = 8'd136; b = 8'd31;  #10 
a = 8'd136; b = 8'd32;  #10 
a = 8'd136; b = 8'd33;  #10 
a = 8'd136; b = 8'd34;  #10 
a = 8'd136; b = 8'd35;  #10 
a = 8'd136; b = 8'd36;  #10 
a = 8'd136; b = 8'd37;  #10 
a = 8'd136; b = 8'd38;  #10 
a = 8'd136; b = 8'd39;  #10 
a = 8'd136; b = 8'd40;  #10 
a = 8'd136; b = 8'd41;  #10 
a = 8'd136; b = 8'd42;  #10 
a = 8'd136; b = 8'd43;  #10 
a = 8'd136; b = 8'd44;  #10 
a = 8'd136; b = 8'd45;  #10 
a = 8'd136; b = 8'd46;  #10 
a = 8'd136; b = 8'd47;  #10 
a = 8'd136; b = 8'd48;  #10 
a = 8'd136; b = 8'd49;  #10 
a = 8'd136; b = 8'd50;  #10 
a = 8'd136; b = 8'd51;  #10 
a = 8'd136; b = 8'd52;  #10 
a = 8'd136; b = 8'd53;  #10 
a = 8'd136; b = 8'd54;  #10 
a = 8'd136; b = 8'd55;  #10 
a = 8'd136; b = 8'd56;  #10 
a = 8'd136; b = 8'd57;  #10 
a = 8'd136; b = 8'd58;  #10 
a = 8'd136; b = 8'd59;  #10 
a = 8'd136; b = 8'd60;  #10 
a = 8'd136; b = 8'd61;  #10 
a = 8'd136; b = 8'd62;  #10 
a = 8'd136; b = 8'd63;  #10 
a = 8'd136; b = 8'd64;  #10 
a = 8'd136; b = 8'd65;  #10 
a = 8'd136; b = 8'd66;  #10 
a = 8'd136; b = 8'd67;  #10 
a = 8'd136; b = 8'd68;  #10 
a = 8'd136; b = 8'd69;  #10 
a = 8'd136; b = 8'd70;  #10 
a = 8'd136; b = 8'd71;  #10 
a = 8'd136; b = 8'd72;  #10 
a = 8'd136; b = 8'd73;  #10 
a = 8'd136; b = 8'd74;  #10 
a = 8'd136; b = 8'd75;  #10 
a = 8'd136; b = 8'd76;  #10 
a = 8'd136; b = 8'd77;  #10 
a = 8'd136; b = 8'd78;  #10 
a = 8'd136; b = 8'd79;  #10 
a = 8'd136; b = 8'd80;  #10 
a = 8'd136; b = 8'd81;  #10 
a = 8'd136; b = 8'd82;  #10 
a = 8'd136; b = 8'd83;  #10 
a = 8'd136; b = 8'd84;  #10 
a = 8'd136; b = 8'd85;  #10 
a = 8'd136; b = 8'd86;  #10 
a = 8'd136; b = 8'd87;  #10 
a = 8'd136; b = 8'd88;  #10 
a = 8'd136; b = 8'd89;  #10 
a = 8'd136; b = 8'd90;  #10 
a = 8'd136; b = 8'd91;  #10 
a = 8'd136; b = 8'd92;  #10 
a = 8'd136; b = 8'd93;  #10 
a = 8'd136; b = 8'd94;  #10 
a = 8'd136; b = 8'd95;  #10 
a = 8'd136; b = 8'd96;  #10 
a = 8'd136; b = 8'd97;  #10 
a = 8'd136; b = 8'd98;  #10 
a = 8'd136; b = 8'd99;  #10 
a = 8'd136; b = 8'd100;  #10 
a = 8'd136; b = 8'd101;  #10 
a = 8'd136; b = 8'd102;  #10 
a = 8'd136; b = 8'd103;  #10 
a = 8'd136; b = 8'd104;  #10 
a = 8'd136; b = 8'd105;  #10 
a = 8'd136; b = 8'd106;  #10 
a = 8'd136; b = 8'd107;  #10 
a = 8'd136; b = 8'd108;  #10 
a = 8'd136; b = 8'd109;  #10 
a = 8'd136; b = 8'd110;  #10 
a = 8'd136; b = 8'd111;  #10 
a = 8'd136; b = 8'd112;  #10 
a = 8'd136; b = 8'd113;  #10 
a = 8'd136; b = 8'd114;  #10 
a = 8'd136; b = 8'd115;  #10 
a = 8'd136; b = 8'd116;  #10 
a = 8'd136; b = 8'd117;  #10 
a = 8'd136; b = 8'd118;  #10 
a = 8'd136; b = 8'd119;  #10 
a = 8'd136; b = 8'd120;  #10 
a = 8'd136; b = 8'd121;  #10 
a = 8'd136; b = 8'd122;  #10 
a = 8'd136; b = 8'd123;  #10 
a = 8'd136; b = 8'd124;  #10 
a = 8'd136; b = 8'd125;  #10 
a = 8'd136; b = 8'd126;  #10 
a = 8'd136; b = 8'd127;  #10 
a = 8'd136; b = 8'd128;  #10 
a = 8'd136; b = 8'd129;  #10 
a = 8'd136; b = 8'd130;  #10 
a = 8'd136; b = 8'd131;  #10 
a = 8'd136; b = 8'd132;  #10 
a = 8'd136; b = 8'd133;  #10 
a = 8'd136; b = 8'd134;  #10 
a = 8'd136; b = 8'd135;  #10 
a = 8'd136; b = 8'd136;  #10 
a = 8'd136; b = 8'd137;  #10 
a = 8'd136; b = 8'd138;  #10 
a = 8'd136; b = 8'd139;  #10 
a = 8'd136; b = 8'd140;  #10 
a = 8'd136; b = 8'd141;  #10 
a = 8'd136; b = 8'd142;  #10 
a = 8'd136; b = 8'd143;  #10 
a = 8'd136; b = 8'd144;  #10 
a = 8'd136; b = 8'd145;  #10 
a = 8'd136; b = 8'd146;  #10 
a = 8'd136; b = 8'd147;  #10 
a = 8'd136; b = 8'd148;  #10 
a = 8'd136; b = 8'd149;  #10 
a = 8'd136; b = 8'd150;  #10 
a = 8'd136; b = 8'd151;  #10 
a = 8'd136; b = 8'd152;  #10 
a = 8'd136; b = 8'd153;  #10 
a = 8'd136; b = 8'd154;  #10 
a = 8'd136; b = 8'd155;  #10 
a = 8'd136; b = 8'd156;  #10 
a = 8'd136; b = 8'd157;  #10 
a = 8'd136; b = 8'd158;  #10 
a = 8'd136; b = 8'd159;  #10 
a = 8'd136; b = 8'd160;  #10 
a = 8'd136; b = 8'd161;  #10 
a = 8'd136; b = 8'd162;  #10 
a = 8'd136; b = 8'd163;  #10 
a = 8'd136; b = 8'd164;  #10 
a = 8'd136; b = 8'd165;  #10 
a = 8'd136; b = 8'd166;  #10 
a = 8'd136; b = 8'd167;  #10 
a = 8'd136; b = 8'd168;  #10 
a = 8'd136; b = 8'd169;  #10 
a = 8'd136; b = 8'd170;  #10 
a = 8'd136; b = 8'd171;  #10 
a = 8'd136; b = 8'd172;  #10 
a = 8'd136; b = 8'd173;  #10 
a = 8'd136; b = 8'd174;  #10 
a = 8'd136; b = 8'd175;  #10 
a = 8'd136; b = 8'd176;  #10 
a = 8'd136; b = 8'd177;  #10 
a = 8'd136; b = 8'd178;  #10 
a = 8'd136; b = 8'd179;  #10 
a = 8'd136; b = 8'd180;  #10 
a = 8'd136; b = 8'd181;  #10 
a = 8'd136; b = 8'd182;  #10 
a = 8'd136; b = 8'd183;  #10 
a = 8'd136; b = 8'd184;  #10 
a = 8'd136; b = 8'd185;  #10 
a = 8'd136; b = 8'd186;  #10 
a = 8'd136; b = 8'd187;  #10 
a = 8'd136; b = 8'd188;  #10 
a = 8'd136; b = 8'd189;  #10 
a = 8'd136; b = 8'd190;  #10 
a = 8'd136; b = 8'd191;  #10 
a = 8'd136; b = 8'd192;  #10 
a = 8'd136; b = 8'd193;  #10 
a = 8'd136; b = 8'd194;  #10 
a = 8'd136; b = 8'd195;  #10 
a = 8'd136; b = 8'd196;  #10 
a = 8'd136; b = 8'd197;  #10 
a = 8'd136; b = 8'd198;  #10 
a = 8'd136; b = 8'd199;  #10 
a = 8'd136; b = 8'd200;  #10 
a = 8'd136; b = 8'd201;  #10 
a = 8'd136; b = 8'd202;  #10 
a = 8'd136; b = 8'd203;  #10 
a = 8'd136; b = 8'd204;  #10 
a = 8'd136; b = 8'd205;  #10 
a = 8'd136; b = 8'd206;  #10 
a = 8'd136; b = 8'd207;  #10 
a = 8'd136; b = 8'd208;  #10 
a = 8'd136; b = 8'd209;  #10 
a = 8'd136; b = 8'd210;  #10 
a = 8'd136; b = 8'd211;  #10 
a = 8'd136; b = 8'd212;  #10 
a = 8'd136; b = 8'd213;  #10 
a = 8'd136; b = 8'd214;  #10 
a = 8'd136; b = 8'd215;  #10 
a = 8'd136; b = 8'd216;  #10 
a = 8'd136; b = 8'd217;  #10 
a = 8'd136; b = 8'd218;  #10 
a = 8'd136; b = 8'd219;  #10 
a = 8'd136; b = 8'd220;  #10 
a = 8'd136; b = 8'd221;  #10 
a = 8'd136; b = 8'd222;  #10 
a = 8'd136; b = 8'd223;  #10 
a = 8'd136; b = 8'd224;  #10 
a = 8'd136; b = 8'd225;  #10 
a = 8'd136; b = 8'd226;  #10 
a = 8'd136; b = 8'd227;  #10 
a = 8'd136; b = 8'd228;  #10 
a = 8'd136; b = 8'd229;  #10 
a = 8'd136; b = 8'd230;  #10 
a = 8'd136; b = 8'd231;  #10 
a = 8'd136; b = 8'd232;  #10 
a = 8'd136; b = 8'd233;  #10 
a = 8'd136; b = 8'd234;  #10 
a = 8'd136; b = 8'd235;  #10 
a = 8'd136; b = 8'd236;  #10 
a = 8'd136; b = 8'd237;  #10 
a = 8'd136; b = 8'd238;  #10 
a = 8'd136; b = 8'd239;  #10 
a = 8'd136; b = 8'd240;  #10 
a = 8'd136; b = 8'd241;  #10 
a = 8'd136; b = 8'd242;  #10 
a = 8'd136; b = 8'd243;  #10 
a = 8'd136; b = 8'd244;  #10 
a = 8'd136; b = 8'd245;  #10 
a = 8'd136; b = 8'd246;  #10 
a = 8'd136; b = 8'd247;  #10 
a = 8'd136; b = 8'd248;  #10 
a = 8'd136; b = 8'd249;  #10 
a = 8'd136; b = 8'd250;  #10 
a = 8'd136; b = 8'd251;  #10 
a = 8'd136; b = 8'd252;  #10 
a = 8'd136; b = 8'd253;  #10 
a = 8'd136; b = 8'd254;  #10 
a = 8'd136; b = 8'd255;  #10 
a = 8'd137; b = 8'd0;  #10 
a = 8'd137; b = 8'd1;  #10 
a = 8'd137; b = 8'd2;  #10 
a = 8'd137; b = 8'd3;  #10 
a = 8'd137; b = 8'd4;  #10 
a = 8'd137; b = 8'd5;  #10 
a = 8'd137; b = 8'd6;  #10 
a = 8'd137; b = 8'd7;  #10 
a = 8'd137; b = 8'd8;  #10 
a = 8'd137; b = 8'd9;  #10 
a = 8'd137; b = 8'd10;  #10 
a = 8'd137; b = 8'd11;  #10 
a = 8'd137; b = 8'd12;  #10 
a = 8'd137; b = 8'd13;  #10 
a = 8'd137; b = 8'd14;  #10 
a = 8'd137; b = 8'd15;  #10 
a = 8'd137; b = 8'd16;  #10 
a = 8'd137; b = 8'd17;  #10 
a = 8'd137; b = 8'd18;  #10 
a = 8'd137; b = 8'd19;  #10 
a = 8'd137; b = 8'd20;  #10 
a = 8'd137; b = 8'd21;  #10 
a = 8'd137; b = 8'd22;  #10 
a = 8'd137; b = 8'd23;  #10 
a = 8'd137; b = 8'd24;  #10 
a = 8'd137; b = 8'd25;  #10 
a = 8'd137; b = 8'd26;  #10 
a = 8'd137; b = 8'd27;  #10 
a = 8'd137; b = 8'd28;  #10 
a = 8'd137; b = 8'd29;  #10 
a = 8'd137; b = 8'd30;  #10 
a = 8'd137; b = 8'd31;  #10 
a = 8'd137; b = 8'd32;  #10 
a = 8'd137; b = 8'd33;  #10 
a = 8'd137; b = 8'd34;  #10 
a = 8'd137; b = 8'd35;  #10 
a = 8'd137; b = 8'd36;  #10 
a = 8'd137; b = 8'd37;  #10 
a = 8'd137; b = 8'd38;  #10 
a = 8'd137; b = 8'd39;  #10 
a = 8'd137; b = 8'd40;  #10 
a = 8'd137; b = 8'd41;  #10 
a = 8'd137; b = 8'd42;  #10 
a = 8'd137; b = 8'd43;  #10 
a = 8'd137; b = 8'd44;  #10 
a = 8'd137; b = 8'd45;  #10 
a = 8'd137; b = 8'd46;  #10 
a = 8'd137; b = 8'd47;  #10 
a = 8'd137; b = 8'd48;  #10 
a = 8'd137; b = 8'd49;  #10 
a = 8'd137; b = 8'd50;  #10 
a = 8'd137; b = 8'd51;  #10 
a = 8'd137; b = 8'd52;  #10 
a = 8'd137; b = 8'd53;  #10 
a = 8'd137; b = 8'd54;  #10 
a = 8'd137; b = 8'd55;  #10 
a = 8'd137; b = 8'd56;  #10 
a = 8'd137; b = 8'd57;  #10 
a = 8'd137; b = 8'd58;  #10 
a = 8'd137; b = 8'd59;  #10 
a = 8'd137; b = 8'd60;  #10 
a = 8'd137; b = 8'd61;  #10 
a = 8'd137; b = 8'd62;  #10 
a = 8'd137; b = 8'd63;  #10 
a = 8'd137; b = 8'd64;  #10 
a = 8'd137; b = 8'd65;  #10 
a = 8'd137; b = 8'd66;  #10 
a = 8'd137; b = 8'd67;  #10 
a = 8'd137; b = 8'd68;  #10 
a = 8'd137; b = 8'd69;  #10 
a = 8'd137; b = 8'd70;  #10 
a = 8'd137; b = 8'd71;  #10 
a = 8'd137; b = 8'd72;  #10 
a = 8'd137; b = 8'd73;  #10 
a = 8'd137; b = 8'd74;  #10 
a = 8'd137; b = 8'd75;  #10 
a = 8'd137; b = 8'd76;  #10 
a = 8'd137; b = 8'd77;  #10 
a = 8'd137; b = 8'd78;  #10 
a = 8'd137; b = 8'd79;  #10 
a = 8'd137; b = 8'd80;  #10 
a = 8'd137; b = 8'd81;  #10 
a = 8'd137; b = 8'd82;  #10 
a = 8'd137; b = 8'd83;  #10 
a = 8'd137; b = 8'd84;  #10 
a = 8'd137; b = 8'd85;  #10 
a = 8'd137; b = 8'd86;  #10 
a = 8'd137; b = 8'd87;  #10 
a = 8'd137; b = 8'd88;  #10 
a = 8'd137; b = 8'd89;  #10 
a = 8'd137; b = 8'd90;  #10 
a = 8'd137; b = 8'd91;  #10 
a = 8'd137; b = 8'd92;  #10 
a = 8'd137; b = 8'd93;  #10 
a = 8'd137; b = 8'd94;  #10 
a = 8'd137; b = 8'd95;  #10 
a = 8'd137; b = 8'd96;  #10 
a = 8'd137; b = 8'd97;  #10 
a = 8'd137; b = 8'd98;  #10 
a = 8'd137; b = 8'd99;  #10 
a = 8'd137; b = 8'd100;  #10 
a = 8'd137; b = 8'd101;  #10 
a = 8'd137; b = 8'd102;  #10 
a = 8'd137; b = 8'd103;  #10 
a = 8'd137; b = 8'd104;  #10 
a = 8'd137; b = 8'd105;  #10 
a = 8'd137; b = 8'd106;  #10 
a = 8'd137; b = 8'd107;  #10 
a = 8'd137; b = 8'd108;  #10 
a = 8'd137; b = 8'd109;  #10 
a = 8'd137; b = 8'd110;  #10 
a = 8'd137; b = 8'd111;  #10 
a = 8'd137; b = 8'd112;  #10 
a = 8'd137; b = 8'd113;  #10 
a = 8'd137; b = 8'd114;  #10 
a = 8'd137; b = 8'd115;  #10 
a = 8'd137; b = 8'd116;  #10 
a = 8'd137; b = 8'd117;  #10 
a = 8'd137; b = 8'd118;  #10 
a = 8'd137; b = 8'd119;  #10 
a = 8'd137; b = 8'd120;  #10 
a = 8'd137; b = 8'd121;  #10 
a = 8'd137; b = 8'd122;  #10 
a = 8'd137; b = 8'd123;  #10 
a = 8'd137; b = 8'd124;  #10 
a = 8'd137; b = 8'd125;  #10 
a = 8'd137; b = 8'd126;  #10 
a = 8'd137; b = 8'd127;  #10 
a = 8'd137; b = 8'd128;  #10 
a = 8'd137; b = 8'd129;  #10 
a = 8'd137; b = 8'd130;  #10 
a = 8'd137; b = 8'd131;  #10 
a = 8'd137; b = 8'd132;  #10 
a = 8'd137; b = 8'd133;  #10 
a = 8'd137; b = 8'd134;  #10 
a = 8'd137; b = 8'd135;  #10 
a = 8'd137; b = 8'd136;  #10 
a = 8'd137; b = 8'd137;  #10 
a = 8'd137; b = 8'd138;  #10 
a = 8'd137; b = 8'd139;  #10 
a = 8'd137; b = 8'd140;  #10 
a = 8'd137; b = 8'd141;  #10 
a = 8'd137; b = 8'd142;  #10 
a = 8'd137; b = 8'd143;  #10 
a = 8'd137; b = 8'd144;  #10 
a = 8'd137; b = 8'd145;  #10 
a = 8'd137; b = 8'd146;  #10 
a = 8'd137; b = 8'd147;  #10 
a = 8'd137; b = 8'd148;  #10 
a = 8'd137; b = 8'd149;  #10 
a = 8'd137; b = 8'd150;  #10 
a = 8'd137; b = 8'd151;  #10 
a = 8'd137; b = 8'd152;  #10 
a = 8'd137; b = 8'd153;  #10 
a = 8'd137; b = 8'd154;  #10 
a = 8'd137; b = 8'd155;  #10 
a = 8'd137; b = 8'd156;  #10 
a = 8'd137; b = 8'd157;  #10 
a = 8'd137; b = 8'd158;  #10 
a = 8'd137; b = 8'd159;  #10 
a = 8'd137; b = 8'd160;  #10 
a = 8'd137; b = 8'd161;  #10 
a = 8'd137; b = 8'd162;  #10 
a = 8'd137; b = 8'd163;  #10 
a = 8'd137; b = 8'd164;  #10 
a = 8'd137; b = 8'd165;  #10 
a = 8'd137; b = 8'd166;  #10 
a = 8'd137; b = 8'd167;  #10 
a = 8'd137; b = 8'd168;  #10 
a = 8'd137; b = 8'd169;  #10 
a = 8'd137; b = 8'd170;  #10 
a = 8'd137; b = 8'd171;  #10 
a = 8'd137; b = 8'd172;  #10 
a = 8'd137; b = 8'd173;  #10 
a = 8'd137; b = 8'd174;  #10 
a = 8'd137; b = 8'd175;  #10 
a = 8'd137; b = 8'd176;  #10 
a = 8'd137; b = 8'd177;  #10 
a = 8'd137; b = 8'd178;  #10 
a = 8'd137; b = 8'd179;  #10 
a = 8'd137; b = 8'd180;  #10 
a = 8'd137; b = 8'd181;  #10 
a = 8'd137; b = 8'd182;  #10 
a = 8'd137; b = 8'd183;  #10 
a = 8'd137; b = 8'd184;  #10 
a = 8'd137; b = 8'd185;  #10 
a = 8'd137; b = 8'd186;  #10 
a = 8'd137; b = 8'd187;  #10 
a = 8'd137; b = 8'd188;  #10 
a = 8'd137; b = 8'd189;  #10 
a = 8'd137; b = 8'd190;  #10 
a = 8'd137; b = 8'd191;  #10 
a = 8'd137; b = 8'd192;  #10 
a = 8'd137; b = 8'd193;  #10 
a = 8'd137; b = 8'd194;  #10 
a = 8'd137; b = 8'd195;  #10 
a = 8'd137; b = 8'd196;  #10 
a = 8'd137; b = 8'd197;  #10 
a = 8'd137; b = 8'd198;  #10 
a = 8'd137; b = 8'd199;  #10 
a = 8'd137; b = 8'd200;  #10 
a = 8'd137; b = 8'd201;  #10 
a = 8'd137; b = 8'd202;  #10 
a = 8'd137; b = 8'd203;  #10 
a = 8'd137; b = 8'd204;  #10 
a = 8'd137; b = 8'd205;  #10 
a = 8'd137; b = 8'd206;  #10 
a = 8'd137; b = 8'd207;  #10 
a = 8'd137; b = 8'd208;  #10 
a = 8'd137; b = 8'd209;  #10 
a = 8'd137; b = 8'd210;  #10 
a = 8'd137; b = 8'd211;  #10 
a = 8'd137; b = 8'd212;  #10 
a = 8'd137; b = 8'd213;  #10 
a = 8'd137; b = 8'd214;  #10 
a = 8'd137; b = 8'd215;  #10 
a = 8'd137; b = 8'd216;  #10 
a = 8'd137; b = 8'd217;  #10 
a = 8'd137; b = 8'd218;  #10 
a = 8'd137; b = 8'd219;  #10 
a = 8'd137; b = 8'd220;  #10 
a = 8'd137; b = 8'd221;  #10 
a = 8'd137; b = 8'd222;  #10 
a = 8'd137; b = 8'd223;  #10 
a = 8'd137; b = 8'd224;  #10 
a = 8'd137; b = 8'd225;  #10 
a = 8'd137; b = 8'd226;  #10 
a = 8'd137; b = 8'd227;  #10 
a = 8'd137; b = 8'd228;  #10 
a = 8'd137; b = 8'd229;  #10 
a = 8'd137; b = 8'd230;  #10 
a = 8'd137; b = 8'd231;  #10 
a = 8'd137; b = 8'd232;  #10 
a = 8'd137; b = 8'd233;  #10 
a = 8'd137; b = 8'd234;  #10 
a = 8'd137; b = 8'd235;  #10 
a = 8'd137; b = 8'd236;  #10 
a = 8'd137; b = 8'd237;  #10 
a = 8'd137; b = 8'd238;  #10 
a = 8'd137; b = 8'd239;  #10 
a = 8'd137; b = 8'd240;  #10 
a = 8'd137; b = 8'd241;  #10 
a = 8'd137; b = 8'd242;  #10 
a = 8'd137; b = 8'd243;  #10 
a = 8'd137; b = 8'd244;  #10 
a = 8'd137; b = 8'd245;  #10 
a = 8'd137; b = 8'd246;  #10 
a = 8'd137; b = 8'd247;  #10 
a = 8'd137; b = 8'd248;  #10 
a = 8'd137; b = 8'd249;  #10 
a = 8'd137; b = 8'd250;  #10 
a = 8'd137; b = 8'd251;  #10 
a = 8'd137; b = 8'd252;  #10 
a = 8'd137; b = 8'd253;  #10 
a = 8'd137; b = 8'd254;  #10 
a = 8'd137; b = 8'd255;  #10 
a = 8'd138; b = 8'd0;  #10 
a = 8'd138; b = 8'd1;  #10 
a = 8'd138; b = 8'd2;  #10 
a = 8'd138; b = 8'd3;  #10 
a = 8'd138; b = 8'd4;  #10 
a = 8'd138; b = 8'd5;  #10 
a = 8'd138; b = 8'd6;  #10 
a = 8'd138; b = 8'd7;  #10 
a = 8'd138; b = 8'd8;  #10 
a = 8'd138; b = 8'd9;  #10 
a = 8'd138; b = 8'd10;  #10 
a = 8'd138; b = 8'd11;  #10 
a = 8'd138; b = 8'd12;  #10 
a = 8'd138; b = 8'd13;  #10 
a = 8'd138; b = 8'd14;  #10 
a = 8'd138; b = 8'd15;  #10 
a = 8'd138; b = 8'd16;  #10 
a = 8'd138; b = 8'd17;  #10 
a = 8'd138; b = 8'd18;  #10 
a = 8'd138; b = 8'd19;  #10 
a = 8'd138; b = 8'd20;  #10 
a = 8'd138; b = 8'd21;  #10 
a = 8'd138; b = 8'd22;  #10 
a = 8'd138; b = 8'd23;  #10 
a = 8'd138; b = 8'd24;  #10 
a = 8'd138; b = 8'd25;  #10 
a = 8'd138; b = 8'd26;  #10 
a = 8'd138; b = 8'd27;  #10 
a = 8'd138; b = 8'd28;  #10 
a = 8'd138; b = 8'd29;  #10 
a = 8'd138; b = 8'd30;  #10 
a = 8'd138; b = 8'd31;  #10 
a = 8'd138; b = 8'd32;  #10 
a = 8'd138; b = 8'd33;  #10 
a = 8'd138; b = 8'd34;  #10 
a = 8'd138; b = 8'd35;  #10 
a = 8'd138; b = 8'd36;  #10 
a = 8'd138; b = 8'd37;  #10 
a = 8'd138; b = 8'd38;  #10 
a = 8'd138; b = 8'd39;  #10 
a = 8'd138; b = 8'd40;  #10 
a = 8'd138; b = 8'd41;  #10 
a = 8'd138; b = 8'd42;  #10 
a = 8'd138; b = 8'd43;  #10 
a = 8'd138; b = 8'd44;  #10 
a = 8'd138; b = 8'd45;  #10 
a = 8'd138; b = 8'd46;  #10 
a = 8'd138; b = 8'd47;  #10 
a = 8'd138; b = 8'd48;  #10 
a = 8'd138; b = 8'd49;  #10 
a = 8'd138; b = 8'd50;  #10 
a = 8'd138; b = 8'd51;  #10 
a = 8'd138; b = 8'd52;  #10 
a = 8'd138; b = 8'd53;  #10 
a = 8'd138; b = 8'd54;  #10 
a = 8'd138; b = 8'd55;  #10 
a = 8'd138; b = 8'd56;  #10 
a = 8'd138; b = 8'd57;  #10 
a = 8'd138; b = 8'd58;  #10 
a = 8'd138; b = 8'd59;  #10 
a = 8'd138; b = 8'd60;  #10 
a = 8'd138; b = 8'd61;  #10 
a = 8'd138; b = 8'd62;  #10 
a = 8'd138; b = 8'd63;  #10 
a = 8'd138; b = 8'd64;  #10 
a = 8'd138; b = 8'd65;  #10 
a = 8'd138; b = 8'd66;  #10 
a = 8'd138; b = 8'd67;  #10 
a = 8'd138; b = 8'd68;  #10 
a = 8'd138; b = 8'd69;  #10 
a = 8'd138; b = 8'd70;  #10 
a = 8'd138; b = 8'd71;  #10 
a = 8'd138; b = 8'd72;  #10 
a = 8'd138; b = 8'd73;  #10 
a = 8'd138; b = 8'd74;  #10 
a = 8'd138; b = 8'd75;  #10 
a = 8'd138; b = 8'd76;  #10 
a = 8'd138; b = 8'd77;  #10 
a = 8'd138; b = 8'd78;  #10 
a = 8'd138; b = 8'd79;  #10 
a = 8'd138; b = 8'd80;  #10 
a = 8'd138; b = 8'd81;  #10 
a = 8'd138; b = 8'd82;  #10 
a = 8'd138; b = 8'd83;  #10 
a = 8'd138; b = 8'd84;  #10 
a = 8'd138; b = 8'd85;  #10 
a = 8'd138; b = 8'd86;  #10 
a = 8'd138; b = 8'd87;  #10 
a = 8'd138; b = 8'd88;  #10 
a = 8'd138; b = 8'd89;  #10 
a = 8'd138; b = 8'd90;  #10 
a = 8'd138; b = 8'd91;  #10 
a = 8'd138; b = 8'd92;  #10 
a = 8'd138; b = 8'd93;  #10 
a = 8'd138; b = 8'd94;  #10 
a = 8'd138; b = 8'd95;  #10 
a = 8'd138; b = 8'd96;  #10 
a = 8'd138; b = 8'd97;  #10 
a = 8'd138; b = 8'd98;  #10 
a = 8'd138; b = 8'd99;  #10 
a = 8'd138; b = 8'd100;  #10 
a = 8'd138; b = 8'd101;  #10 
a = 8'd138; b = 8'd102;  #10 
a = 8'd138; b = 8'd103;  #10 
a = 8'd138; b = 8'd104;  #10 
a = 8'd138; b = 8'd105;  #10 
a = 8'd138; b = 8'd106;  #10 
a = 8'd138; b = 8'd107;  #10 
a = 8'd138; b = 8'd108;  #10 
a = 8'd138; b = 8'd109;  #10 
a = 8'd138; b = 8'd110;  #10 
a = 8'd138; b = 8'd111;  #10 
a = 8'd138; b = 8'd112;  #10 
a = 8'd138; b = 8'd113;  #10 
a = 8'd138; b = 8'd114;  #10 
a = 8'd138; b = 8'd115;  #10 
a = 8'd138; b = 8'd116;  #10 
a = 8'd138; b = 8'd117;  #10 
a = 8'd138; b = 8'd118;  #10 
a = 8'd138; b = 8'd119;  #10 
a = 8'd138; b = 8'd120;  #10 
a = 8'd138; b = 8'd121;  #10 
a = 8'd138; b = 8'd122;  #10 
a = 8'd138; b = 8'd123;  #10 
a = 8'd138; b = 8'd124;  #10 
a = 8'd138; b = 8'd125;  #10 
a = 8'd138; b = 8'd126;  #10 
a = 8'd138; b = 8'd127;  #10 
a = 8'd138; b = 8'd128;  #10 
a = 8'd138; b = 8'd129;  #10 
a = 8'd138; b = 8'd130;  #10 
a = 8'd138; b = 8'd131;  #10 
a = 8'd138; b = 8'd132;  #10 
a = 8'd138; b = 8'd133;  #10 
a = 8'd138; b = 8'd134;  #10 
a = 8'd138; b = 8'd135;  #10 
a = 8'd138; b = 8'd136;  #10 
a = 8'd138; b = 8'd137;  #10 
a = 8'd138; b = 8'd138;  #10 
a = 8'd138; b = 8'd139;  #10 
a = 8'd138; b = 8'd140;  #10 
a = 8'd138; b = 8'd141;  #10 
a = 8'd138; b = 8'd142;  #10 
a = 8'd138; b = 8'd143;  #10 
a = 8'd138; b = 8'd144;  #10 
a = 8'd138; b = 8'd145;  #10 
a = 8'd138; b = 8'd146;  #10 
a = 8'd138; b = 8'd147;  #10 
a = 8'd138; b = 8'd148;  #10 
a = 8'd138; b = 8'd149;  #10 
a = 8'd138; b = 8'd150;  #10 
a = 8'd138; b = 8'd151;  #10 
a = 8'd138; b = 8'd152;  #10 
a = 8'd138; b = 8'd153;  #10 
a = 8'd138; b = 8'd154;  #10 
a = 8'd138; b = 8'd155;  #10 
a = 8'd138; b = 8'd156;  #10 
a = 8'd138; b = 8'd157;  #10 
a = 8'd138; b = 8'd158;  #10 
a = 8'd138; b = 8'd159;  #10 
a = 8'd138; b = 8'd160;  #10 
a = 8'd138; b = 8'd161;  #10 
a = 8'd138; b = 8'd162;  #10 
a = 8'd138; b = 8'd163;  #10 
a = 8'd138; b = 8'd164;  #10 
a = 8'd138; b = 8'd165;  #10 
a = 8'd138; b = 8'd166;  #10 
a = 8'd138; b = 8'd167;  #10 
a = 8'd138; b = 8'd168;  #10 
a = 8'd138; b = 8'd169;  #10 
a = 8'd138; b = 8'd170;  #10 
a = 8'd138; b = 8'd171;  #10 
a = 8'd138; b = 8'd172;  #10 
a = 8'd138; b = 8'd173;  #10 
a = 8'd138; b = 8'd174;  #10 
a = 8'd138; b = 8'd175;  #10 
a = 8'd138; b = 8'd176;  #10 
a = 8'd138; b = 8'd177;  #10 
a = 8'd138; b = 8'd178;  #10 
a = 8'd138; b = 8'd179;  #10 
a = 8'd138; b = 8'd180;  #10 
a = 8'd138; b = 8'd181;  #10 
a = 8'd138; b = 8'd182;  #10 
a = 8'd138; b = 8'd183;  #10 
a = 8'd138; b = 8'd184;  #10 
a = 8'd138; b = 8'd185;  #10 
a = 8'd138; b = 8'd186;  #10 
a = 8'd138; b = 8'd187;  #10 
a = 8'd138; b = 8'd188;  #10 
a = 8'd138; b = 8'd189;  #10 
a = 8'd138; b = 8'd190;  #10 
a = 8'd138; b = 8'd191;  #10 
a = 8'd138; b = 8'd192;  #10 
a = 8'd138; b = 8'd193;  #10 
a = 8'd138; b = 8'd194;  #10 
a = 8'd138; b = 8'd195;  #10 
a = 8'd138; b = 8'd196;  #10 
a = 8'd138; b = 8'd197;  #10 
a = 8'd138; b = 8'd198;  #10 
a = 8'd138; b = 8'd199;  #10 
a = 8'd138; b = 8'd200;  #10 
a = 8'd138; b = 8'd201;  #10 
a = 8'd138; b = 8'd202;  #10 
a = 8'd138; b = 8'd203;  #10 
a = 8'd138; b = 8'd204;  #10 
a = 8'd138; b = 8'd205;  #10 
a = 8'd138; b = 8'd206;  #10 
a = 8'd138; b = 8'd207;  #10 
a = 8'd138; b = 8'd208;  #10 
a = 8'd138; b = 8'd209;  #10 
a = 8'd138; b = 8'd210;  #10 
a = 8'd138; b = 8'd211;  #10 
a = 8'd138; b = 8'd212;  #10 
a = 8'd138; b = 8'd213;  #10 
a = 8'd138; b = 8'd214;  #10 
a = 8'd138; b = 8'd215;  #10 
a = 8'd138; b = 8'd216;  #10 
a = 8'd138; b = 8'd217;  #10 
a = 8'd138; b = 8'd218;  #10 
a = 8'd138; b = 8'd219;  #10 
a = 8'd138; b = 8'd220;  #10 
a = 8'd138; b = 8'd221;  #10 
a = 8'd138; b = 8'd222;  #10 
a = 8'd138; b = 8'd223;  #10 
a = 8'd138; b = 8'd224;  #10 
a = 8'd138; b = 8'd225;  #10 
a = 8'd138; b = 8'd226;  #10 
a = 8'd138; b = 8'd227;  #10 
a = 8'd138; b = 8'd228;  #10 
a = 8'd138; b = 8'd229;  #10 
a = 8'd138; b = 8'd230;  #10 
a = 8'd138; b = 8'd231;  #10 
a = 8'd138; b = 8'd232;  #10 
a = 8'd138; b = 8'd233;  #10 
a = 8'd138; b = 8'd234;  #10 
a = 8'd138; b = 8'd235;  #10 
a = 8'd138; b = 8'd236;  #10 
a = 8'd138; b = 8'd237;  #10 
a = 8'd138; b = 8'd238;  #10 
a = 8'd138; b = 8'd239;  #10 
a = 8'd138; b = 8'd240;  #10 
a = 8'd138; b = 8'd241;  #10 
a = 8'd138; b = 8'd242;  #10 
a = 8'd138; b = 8'd243;  #10 
a = 8'd138; b = 8'd244;  #10 
a = 8'd138; b = 8'd245;  #10 
a = 8'd138; b = 8'd246;  #10 
a = 8'd138; b = 8'd247;  #10 
a = 8'd138; b = 8'd248;  #10 
a = 8'd138; b = 8'd249;  #10 
a = 8'd138; b = 8'd250;  #10 
a = 8'd138; b = 8'd251;  #10 
a = 8'd138; b = 8'd252;  #10 
a = 8'd138; b = 8'd253;  #10 
a = 8'd138; b = 8'd254;  #10 
a = 8'd138; b = 8'd255;  #10 
a = 8'd139; b = 8'd0;  #10 
a = 8'd139; b = 8'd1;  #10 
a = 8'd139; b = 8'd2;  #10 
a = 8'd139; b = 8'd3;  #10 
a = 8'd139; b = 8'd4;  #10 
a = 8'd139; b = 8'd5;  #10 
a = 8'd139; b = 8'd6;  #10 
a = 8'd139; b = 8'd7;  #10 
a = 8'd139; b = 8'd8;  #10 
a = 8'd139; b = 8'd9;  #10 
a = 8'd139; b = 8'd10;  #10 
a = 8'd139; b = 8'd11;  #10 
a = 8'd139; b = 8'd12;  #10 
a = 8'd139; b = 8'd13;  #10 
a = 8'd139; b = 8'd14;  #10 
a = 8'd139; b = 8'd15;  #10 
a = 8'd139; b = 8'd16;  #10 
a = 8'd139; b = 8'd17;  #10 
a = 8'd139; b = 8'd18;  #10 
a = 8'd139; b = 8'd19;  #10 
a = 8'd139; b = 8'd20;  #10 
a = 8'd139; b = 8'd21;  #10 
a = 8'd139; b = 8'd22;  #10 
a = 8'd139; b = 8'd23;  #10 
a = 8'd139; b = 8'd24;  #10 
a = 8'd139; b = 8'd25;  #10 
a = 8'd139; b = 8'd26;  #10 
a = 8'd139; b = 8'd27;  #10 
a = 8'd139; b = 8'd28;  #10 
a = 8'd139; b = 8'd29;  #10 
a = 8'd139; b = 8'd30;  #10 
a = 8'd139; b = 8'd31;  #10 
a = 8'd139; b = 8'd32;  #10 
a = 8'd139; b = 8'd33;  #10 
a = 8'd139; b = 8'd34;  #10 
a = 8'd139; b = 8'd35;  #10 
a = 8'd139; b = 8'd36;  #10 
a = 8'd139; b = 8'd37;  #10 
a = 8'd139; b = 8'd38;  #10 
a = 8'd139; b = 8'd39;  #10 
a = 8'd139; b = 8'd40;  #10 
a = 8'd139; b = 8'd41;  #10 
a = 8'd139; b = 8'd42;  #10 
a = 8'd139; b = 8'd43;  #10 
a = 8'd139; b = 8'd44;  #10 
a = 8'd139; b = 8'd45;  #10 
a = 8'd139; b = 8'd46;  #10 
a = 8'd139; b = 8'd47;  #10 
a = 8'd139; b = 8'd48;  #10 
a = 8'd139; b = 8'd49;  #10 
a = 8'd139; b = 8'd50;  #10 
a = 8'd139; b = 8'd51;  #10 
a = 8'd139; b = 8'd52;  #10 
a = 8'd139; b = 8'd53;  #10 
a = 8'd139; b = 8'd54;  #10 
a = 8'd139; b = 8'd55;  #10 
a = 8'd139; b = 8'd56;  #10 
a = 8'd139; b = 8'd57;  #10 
a = 8'd139; b = 8'd58;  #10 
a = 8'd139; b = 8'd59;  #10 
a = 8'd139; b = 8'd60;  #10 
a = 8'd139; b = 8'd61;  #10 
a = 8'd139; b = 8'd62;  #10 
a = 8'd139; b = 8'd63;  #10 
a = 8'd139; b = 8'd64;  #10 
a = 8'd139; b = 8'd65;  #10 
a = 8'd139; b = 8'd66;  #10 
a = 8'd139; b = 8'd67;  #10 
a = 8'd139; b = 8'd68;  #10 
a = 8'd139; b = 8'd69;  #10 
a = 8'd139; b = 8'd70;  #10 
a = 8'd139; b = 8'd71;  #10 
a = 8'd139; b = 8'd72;  #10 
a = 8'd139; b = 8'd73;  #10 
a = 8'd139; b = 8'd74;  #10 
a = 8'd139; b = 8'd75;  #10 
a = 8'd139; b = 8'd76;  #10 
a = 8'd139; b = 8'd77;  #10 
a = 8'd139; b = 8'd78;  #10 
a = 8'd139; b = 8'd79;  #10 
a = 8'd139; b = 8'd80;  #10 
a = 8'd139; b = 8'd81;  #10 
a = 8'd139; b = 8'd82;  #10 
a = 8'd139; b = 8'd83;  #10 
a = 8'd139; b = 8'd84;  #10 
a = 8'd139; b = 8'd85;  #10 
a = 8'd139; b = 8'd86;  #10 
a = 8'd139; b = 8'd87;  #10 
a = 8'd139; b = 8'd88;  #10 
a = 8'd139; b = 8'd89;  #10 
a = 8'd139; b = 8'd90;  #10 
a = 8'd139; b = 8'd91;  #10 
a = 8'd139; b = 8'd92;  #10 
a = 8'd139; b = 8'd93;  #10 
a = 8'd139; b = 8'd94;  #10 
a = 8'd139; b = 8'd95;  #10 
a = 8'd139; b = 8'd96;  #10 
a = 8'd139; b = 8'd97;  #10 
a = 8'd139; b = 8'd98;  #10 
a = 8'd139; b = 8'd99;  #10 
a = 8'd139; b = 8'd100;  #10 
a = 8'd139; b = 8'd101;  #10 
a = 8'd139; b = 8'd102;  #10 
a = 8'd139; b = 8'd103;  #10 
a = 8'd139; b = 8'd104;  #10 
a = 8'd139; b = 8'd105;  #10 
a = 8'd139; b = 8'd106;  #10 
a = 8'd139; b = 8'd107;  #10 
a = 8'd139; b = 8'd108;  #10 
a = 8'd139; b = 8'd109;  #10 
a = 8'd139; b = 8'd110;  #10 
a = 8'd139; b = 8'd111;  #10 
a = 8'd139; b = 8'd112;  #10 
a = 8'd139; b = 8'd113;  #10 
a = 8'd139; b = 8'd114;  #10 
a = 8'd139; b = 8'd115;  #10 
a = 8'd139; b = 8'd116;  #10 
a = 8'd139; b = 8'd117;  #10 
a = 8'd139; b = 8'd118;  #10 
a = 8'd139; b = 8'd119;  #10 
a = 8'd139; b = 8'd120;  #10 
a = 8'd139; b = 8'd121;  #10 
a = 8'd139; b = 8'd122;  #10 
a = 8'd139; b = 8'd123;  #10 
a = 8'd139; b = 8'd124;  #10 
a = 8'd139; b = 8'd125;  #10 
a = 8'd139; b = 8'd126;  #10 
a = 8'd139; b = 8'd127;  #10 
a = 8'd139; b = 8'd128;  #10 
a = 8'd139; b = 8'd129;  #10 
a = 8'd139; b = 8'd130;  #10 
a = 8'd139; b = 8'd131;  #10 
a = 8'd139; b = 8'd132;  #10 
a = 8'd139; b = 8'd133;  #10 
a = 8'd139; b = 8'd134;  #10 
a = 8'd139; b = 8'd135;  #10 
a = 8'd139; b = 8'd136;  #10 
a = 8'd139; b = 8'd137;  #10 
a = 8'd139; b = 8'd138;  #10 
a = 8'd139; b = 8'd139;  #10 
a = 8'd139; b = 8'd140;  #10 
a = 8'd139; b = 8'd141;  #10 
a = 8'd139; b = 8'd142;  #10 
a = 8'd139; b = 8'd143;  #10 
a = 8'd139; b = 8'd144;  #10 
a = 8'd139; b = 8'd145;  #10 
a = 8'd139; b = 8'd146;  #10 
a = 8'd139; b = 8'd147;  #10 
a = 8'd139; b = 8'd148;  #10 
a = 8'd139; b = 8'd149;  #10 
a = 8'd139; b = 8'd150;  #10 
a = 8'd139; b = 8'd151;  #10 
a = 8'd139; b = 8'd152;  #10 
a = 8'd139; b = 8'd153;  #10 
a = 8'd139; b = 8'd154;  #10 
a = 8'd139; b = 8'd155;  #10 
a = 8'd139; b = 8'd156;  #10 
a = 8'd139; b = 8'd157;  #10 
a = 8'd139; b = 8'd158;  #10 
a = 8'd139; b = 8'd159;  #10 
a = 8'd139; b = 8'd160;  #10 
a = 8'd139; b = 8'd161;  #10 
a = 8'd139; b = 8'd162;  #10 
a = 8'd139; b = 8'd163;  #10 
a = 8'd139; b = 8'd164;  #10 
a = 8'd139; b = 8'd165;  #10 
a = 8'd139; b = 8'd166;  #10 
a = 8'd139; b = 8'd167;  #10 
a = 8'd139; b = 8'd168;  #10 
a = 8'd139; b = 8'd169;  #10 
a = 8'd139; b = 8'd170;  #10 
a = 8'd139; b = 8'd171;  #10 
a = 8'd139; b = 8'd172;  #10 
a = 8'd139; b = 8'd173;  #10 
a = 8'd139; b = 8'd174;  #10 
a = 8'd139; b = 8'd175;  #10 
a = 8'd139; b = 8'd176;  #10 
a = 8'd139; b = 8'd177;  #10 
a = 8'd139; b = 8'd178;  #10 
a = 8'd139; b = 8'd179;  #10 
a = 8'd139; b = 8'd180;  #10 
a = 8'd139; b = 8'd181;  #10 
a = 8'd139; b = 8'd182;  #10 
a = 8'd139; b = 8'd183;  #10 
a = 8'd139; b = 8'd184;  #10 
a = 8'd139; b = 8'd185;  #10 
a = 8'd139; b = 8'd186;  #10 
a = 8'd139; b = 8'd187;  #10 
a = 8'd139; b = 8'd188;  #10 
a = 8'd139; b = 8'd189;  #10 
a = 8'd139; b = 8'd190;  #10 
a = 8'd139; b = 8'd191;  #10 
a = 8'd139; b = 8'd192;  #10 
a = 8'd139; b = 8'd193;  #10 
a = 8'd139; b = 8'd194;  #10 
a = 8'd139; b = 8'd195;  #10 
a = 8'd139; b = 8'd196;  #10 
a = 8'd139; b = 8'd197;  #10 
a = 8'd139; b = 8'd198;  #10 
a = 8'd139; b = 8'd199;  #10 
a = 8'd139; b = 8'd200;  #10 
a = 8'd139; b = 8'd201;  #10 
a = 8'd139; b = 8'd202;  #10 
a = 8'd139; b = 8'd203;  #10 
a = 8'd139; b = 8'd204;  #10 
a = 8'd139; b = 8'd205;  #10 
a = 8'd139; b = 8'd206;  #10 
a = 8'd139; b = 8'd207;  #10 
a = 8'd139; b = 8'd208;  #10 
a = 8'd139; b = 8'd209;  #10 
a = 8'd139; b = 8'd210;  #10 
a = 8'd139; b = 8'd211;  #10 
a = 8'd139; b = 8'd212;  #10 
a = 8'd139; b = 8'd213;  #10 
a = 8'd139; b = 8'd214;  #10 
a = 8'd139; b = 8'd215;  #10 
a = 8'd139; b = 8'd216;  #10 
a = 8'd139; b = 8'd217;  #10 
a = 8'd139; b = 8'd218;  #10 
a = 8'd139; b = 8'd219;  #10 
a = 8'd139; b = 8'd220;  #10 
a = 8'd139; b = 8'd221;  #10 
a = 8'd139; b = 8'd222;  #10 
a = 8'd139; b = 8'd223;  #10 
a = 8'd139; b = 8'd224;  #10 
a = 8'd139; b = 8'd225;  #10 
a = 8'd139; b = 8'd226;  #10 
a = 8'd139; b = 8'd227;  #10 
a = 8'd139; b = 8'd228;  #10 
a = 8'd139; b = 8'd229;  #10 
a = 8'd139; b = 8'd230;  #10 
a = 8'd139; b = 8'd231;  #10 
a = 8'd139; b = 8'd232;  #10 
a = 8'd139; b = 8'd233;  #10 
a = 8'd139; b = 8'd234;  #10 
a = 8'd139; b = 8'd235;  #10 
a = 8'd139; b = 8'd236;  #10 
a = 8'd139; b = 8'd237;  #10 
a = 8'd139; b = 8'd238;  #10 
a = 8'd139; b = 8'd239;  #10 
a = 8'd139; b = 8'd240;  #10 
a = 8'd139; b = 8'd241;  #10 
a = 8'd139; b = 8'd242;  #10 
a = 8'd139; b = 8'd243;  #10 
a = 8'd139; b = 8'd244;  #10 
a = 8'd139; b = 8'd245;  #10 
a = 8'd139; b = 8'd246;  #10 
a = 8'd139; b = 8'd247;  #10 
a = 8'd139; b = 8'd248;  #10 
a = 8'd139; b = 8'd249;  #10 
a = 8'd139; b = 8'd250;  #10 
a = 8'd139; b = 8'd251;  #10 
a = 8'd139; b = 8'd252;  #10 
a = 8'd139; b = 8'd253;  #10 
a = 8'd139; b = 8'd254;  #10 
a = 8'd139; b = 8'd255;  #10 
a = 8'd140; b = 8'd0;  #10 
a = 8'd140; b = 8'd1;  #10 
a = 8'd140; b = 8'd2;  #10 
a = 8'd140; b = 8'd3;  #10 
a = 8'd140; b = 8'd4;  #10 
a = 8'd140; b = 8'd5;  #10 
a = 8'd140; b = 8'd6;  #10 
a = 8'd140; b = 8'd7;  #10 
a = 8'd140; b = 8'd8;  #10 
a = 8'd140; b = 8'd9;  #10 
a = 8'd140; b = 8'd10;  #10 
a = 8'd140; b = 8'd11;  #10 
a = 8'd140; b = 8'd12;  #10 
a = 8'd140; b = 8'd13;  #10 
a = 8'd140; b = 8'd14;  #10 
a = 8'd140; b = 8'd15;  #10 
a = 8'd140; b = 8'd16;  #10 
a = 8'd140; b = 8'd17;  #10 
a = 8'd140; b = 8'd18;  #10 
a = 8'd140; b = 8'd19;  #10 
a = 8'd140; b = 8'd20;  #10 
a = 8'd140; b = 8'd21;  #10 
a = 8'd140; b = 8'd22;  #10 
a = 8'd140; b = 8'd23;  #10 
a = 8'd140; b = 8'd24;  #10 
a = 8'd140; b = 8'd25;  #10 
a = 8'd140; b = 8'd26;  #10 
a = 8'd140; b = 8'd27;  #10 
a = 8'd140; b = 8'd28;  #10 
a = 8'd140; b = 8'd29;  #10 
a = 8'd140; b = 8'd30;  #10 
a = 8'd140; b = 8'd31;  #10 
a = 8'd140; b = 8'd32;  #10 
a = 8'd140; b = 8'd33;  #10 
a = 8'd140; b = 8'd34;  #10 
a = 8'd140; b = 8'd35;  #10 
a = 8'd140; b = 8'd36;  #10 
a = 8'd140; b = 8'd37;  #10 
a = 8'd140; b = 8'd38;  #10 
a = 8'd140; b = 8'd39;  #10 
a = 8'd140; b = 8'd40;  #10 
a = 8'd140; b = 8'd41;  #10 
a = 8'd140; b = 8'd42;  #10 
a = 8'd140; b = 8'd43;  #10 
a = 8'd140; b = 8'd44;  #10 
a = 8'd140; b = 8'd45;  #10 
a = 8'd140; b = 8'd46;  #10 
a = 8'd140; b = 8'd47;  #10 
a = 8'd140; b = 8'd48;  #10 
a = 8'd140; b = 8'd49;  #10 
a = 8'd140; b = 8'd50;  #10 
a = 8'd140; b = 8'd51;  #10 
a = 8'd140; b = 8'd52;  #10 
a = 8'd140; b = 8'd53;  #10 
a = 8'd140; b = 8'd54;  #10 
a = 8'd140; b = 8'd55;  #10 
a = 8'd140; b = 8'd56;  #10 
a = 8'd140; b = 8'd57;  #10 
a = 8'd140; b = 8'd58;  #10 
a = 8'd140; b = 8'd59;  #10 
a = 8'd140; b = 8'd60;  #10 
a = 8'd140; b = 8'd61;  #10 
a = 8'd140; b = 8'd62;  #10 
a = 8'd140; b = 8'd63;  #10 
a = 8'd140; b = 8'd64;  #10 
a = 8'd140; b = 8'd65;  #10 
a = 8'd140; b = 8'd66;  #10 
a = 8'd140; b = 8'd67;  #10 
a = 8'd140; b = 8'd68;  #10 
a = 8'd140; b = 8'd69;  #10 
a = 8'd140; b = 8'd70;  #10 
a = 8'd140; b = 8'd71;  #10 
a = 8'd140; b = 8'd72;  #10 
a = 8'd140; b = 8'd73;  #10 
a = 8'd140; b = 8'd74;  #10 
a = 8'd140; b = 8'd75;  #10 
a = 8'd140; b = 8'd76;  #10 
a = 8'd140; b = 8'd77;  #10 
a = 8'd140; b = 8'd78;  #10 
a = 8'd140; b = 8'd79;  #10 
a = 8'd140; b = 8'd80;  #10 
a = 8'd140; b = 8'd81;  #10 
a = 8'd140; b = 8'd82;  #10 
a = 8'd140; b = 8'd83;  #10 
a = 8'd140; b = 8'd84;  #10 
a = 8'd140; b = 8'd85;  #10 
a = 8'd140; b = 8'd86;  #10 
a = 8'd140; b = 8'd87;  #10 
a = 8'd140; b = 8'd88;  #10 
a = 8'd140; b = 8'd89;  #10 
a = 8'd140; b = 8'd90;  #10 
a = 8'd140; b = 8'd91;  #10 
a = 8'd140; b = 8'd92;  #10 
a = 8'd140; b = 8'd93;  #10 
a = 8'd140; b = 8'd94;  #10 
a = 8'd140; b = 8'd95;  #10 
a = 8'd140; b = 8'd96;  #10 
a = 8'd140; b = 8'd97;  #10 
a = 8'd140; b = 8'd98;  #10 
a = 8'd140; b = 8'd99;  #10 
a = 8'd140; b = 8'd100;  #10 
a = 8'd140; b = 8'd101;  #10 
a = 8'd140; b = 8'd102;  #10 
a = 8'd140; b = 8'd103;  #10 
a = 8'd140; b = 8'd104;  #10 
a = 8'd140; b = 8'd105;  #10 
a = 8'd140; b = 8'd106;  #10 
a = 8'd140; b = 8'd107;  #10 
a = 8'd140; b = 8'd108;  #10 
a = 8'd140; b = 8'd109;  #10 
a = 8'd140; b = 8'd110;  #10 
a = 8'd140; b = 8'd111;  #10 
a = 8'd140; b = 8'd112;  #10 
a = 8'd140; b = 8'd113;  #10 
a = 8'd140; b = 8'd114;  #10 
a = 8'd140; b = 8'd115;  #10 
a = 8'd140; b = 8'd116;  #10 
a = 8'd140; b = 8'd117;  #10 
a = 8'd140; b = 8'd118;  #10 
a = 8'd140; b = 8'd119;  #10 
a = 8'd140; b = 8'd120;  #10 
a = 8'd140; b = 8'd121;  #10 
a = 8'd140; b = 8'd122;  #10 
a = 8'd140; b = 8'd123;  #10 
a = 8'd140; b = 8'd124;  #10 
a = 8'd140; b = 8'd125;  #10 
a = 8'd140; b = 8'd126;  #10 
a = 8'd140; b = 8'd127;  #10 
a = 8'd140; b = 8'd128;  #10 
a = 8'd140; b = 8'd129;  #10 
a = 8'd140; b = 8'd130;  #10 
a = 8'd140; b = 8'd131;  #10 
a = 8'd140; b = 8'd132;  #10 
a = 8'd140; b = 8'd133;  #10 
a = 8'd140; b = 8'd134;  #10 
a = 8'd140; b = 8'd135;  #10 
a = 8'd140; b = 8'd136;  #10 
a = 8'd140; b = 8'd137;  #10 
a = 8'd140; b = 8'd138;  #10 
a = 8'd140; b = 8'd139;  #10 
a = 8'd140; b = 8'd140;  #10 
a = 8'd140; b = 8'd141;  #10 
a = 8'd140; b = 8'd142;  #10 
a = 8'd140; b = 8'd143;  #10 
a = 8'd140; b = 8'd144;  #10 
a = 8'd140; b = 8'd145;  #10 
a = 8'd140; b = 8'd146;  #10 
a = 8'd140; b = 8'd147;  #10 
a = 8'd140; b = 8'd148;  #10 
a = 8'd140; b = 8'd149;  #10 
a = 8'd140; b = 8'd150;  #10 
a = 8'd140; b = 8'd151;  #10 
a = 8'd140; b = 8'd152;  #10 
a = 8'd140; b = 8'd153;  #10 
a = 8'd140; b = 8'd154;  #10 
a = 8'd140; b = 8'd155;  #10 
a = 8'd140; b = 8'd156;  #10 
a = 8'd140; b = 8'd157;  #10 
a = 8'd140; b = 8'd158;  #10 
a = 8'd140; b = 8'd159;  #10 
a = 8'd140; b = 8'd160;  #10 
a = 8'd140; b = 8'd161;  #10 
a = 8'd140; b = 8'd162;  #10 
a = 8'd140; b = 8'd163;  #10 
a = 8'd140; b = 8'd164;  #10 
a = 8'd140; b = 8'd165;  #10 
a = 8'd140; b = 8'd166;  #10 
a = 8'd140; b = 8'd167;  #10 
a = 8'd140; b = 8'd168;  #10 
a = 8'd140; b = 8'd169;  #10 
a = 8'd140; b = 8'd170;  #10 
a = 8'd140; b = 8'd171;  #10 
a = 8'd140; b = 8'd172;  #10 
a = 8'd140; b = 8'd173;  #10 
a = 8'd140; b = 8'd174;  #10 
a = 8'd140; b = 8'd175;  #10 
a = 8'd140; b = 8'd176;  #10 
a = 8'd140; b = 8'd177;  #10 
a = 8'd140; b = 8'd178;  #10 
a = 8'd140; b = 8'd179;  #10 
a = 8'd140; b = 8'd180;  #10 
a = 8'd140; b = 8'd181;  #10 
a = 8'd140; b = 8'd182;  #10 
a = 8'd140; b = 8'd183;  #10 
a = 8'd140; b = 8'd184;  #10 
a = 8'd140; b = 8'd185;  #10 
a = 8'd140; b = 8'd186;  #10 
a = 8'd140; b = 8'd187;  #10 
a = 8'd140; b = 8'd188;  #10 
a = 8'd140; b = 8'd189;  #10 
a = 8'd140; b = 8'd190;  #10 
a = 8'd140; b = 8'd191;  #10 
a = 8'd140; b = 8'd192;  #10 
a = 8'd140; b = 8'd193;  #10 
a = 8'd140; b = 8'd194;  #10 
a = 8'd140; b = 8'd195;  #10 
a = 8'd140; b = 8'd196;  #10 
a = 8'd140; b = 8'd197;  #10 
a = 8'd140; b = 8'd198;  #10 
a = 8'd140; b = 8'd199;  #10 
a = 8'd140; b = 8'd200;  #10 
a = 8'd140; b = 8'd201;  #10 
a = 8'd140; b = 8'd202;  #10 
a = 8'd140; b = 8'd203;  #10 
a = 8'd140; b = 8'd204;  #10 
a = 8'd140; b = 8'd205;  #10 
a = 8'd140; b = 8'd206;  #10 
a = 8'd140; b = 8'd207;  #10 
a = 8'd140; b = 8'd208;  #10 
a = 8'd140; b = 8'd209;  #10 
a = 8'd140; b = 8'd210;  #10 
a = 8'd140; b = 8'd211;  #10 
a = 8'd140; b = 8'd212;  #10 
a = 8'd140; b = 8'd213;  #10 
a = 8'd140; b = 8'd214;  #10 
a = 8'd140; b = 8'd215;  #10 
a = 8'd140; b = 8'd216;  #10 
a = 8'd140; b = 8'd217;  #10 
a = 8'd140; b = 8'd218;  #10 
a = 8'd140; b = 8'd219;  #10 
a = 8'd140; b = 8'd220;  #10 
a = 8'd140; b = 8'd221;  #10 
a = 8'd140; b = 8'd222;  #10 
a = 8'd140; b = 8'd223;  #10 
a = 8'd140; b = 8'd224;  #10 
a = 8'd140; b = 8'd225;  #10 
a = 8'd140; b = 8'd226;  #10 
a = 8'd140; b = 8'd227;  #10 
a = 8'd140; b = 8'd228;  #10 
a = 8'd140; b = 8'd229;  #10 
a = 8'd140; b = 8'd230;  #10 
a = 8'd140; b = 8'd231;  #10 
a = 8'd140; b = 8'd232;  #10 
a = 8'd140; b = 8'd233;  #10 
a = 8'd140; b = 8'd234;  #10 
a = 8'd140; b = 8'd235;  #10 
a = 8'd140; b = 8'd236;  #10 
a = 8'd140; b = 8'd237;  #10 
a = 8'd140; b = 8'd238;  #10 
a = 8'd140; b = 8'd239;  #10 
a = 8'd140; b = 8'd240;  #10 
a = 8'd140; b = 8'd241;  #10 
a = 8'd140; b = 8'd242;  #10 
a = 8'd140; b = 8'd243;  #10 
a = 8'd140; b = 8'd244;  #10 
a = 8'd140; b = 8'd245;  #10 
a = 8'd140; b = 8'd246;  #10 
a = 8'd140; b = 8'd247;  #10 
a = 8'd140; b = 8'd248;  #10 
a = 8'd140; b = 8'd249;  #10 
a = 8'd140; b = 8'd250;  #10 
a = 8'd140; b = 8'd251;  #10 
a = 8'd140; b = 8'd252;  #10 
a = 8'd140; b = 8'd253;  #10 
a = 8'd140; b = 8'd254;  #10 
a = 8'd140; b = 8'd255;  #10 
a = 8'd141; b = 8'd0;  #10 
a = 8'd141; b = 8'd1;  #10 
a = 8'd141; b = 8'd2;  #10 
a = 8'd141; b = 8'd3;  #10 
a = 8'd141; b = 8'd4;  #10 
a = 8'd141; b = 8'd5;  #10 
a = 8'd141; b = 8'd6;  #10 
a = 8'd141; b = 8'd7;  #10 
a = 8'd141; b = 8'd8;  #10 
a = 8'd141; b = 8'd9;  #10 
a = 8'd141; b = 8'd10;  #10 
a = 8'd141; b = 8'd11;  #10 
a = 8'd141; b = 8'd12;  #10 
a = 8'd141; b = 8'd13;  #10 
a = 8'd141; b = 8'd14;  #10 
a = 8'd141; b = 8'd15;  #10 
a = 8'd141; b = 8'd16;  #10 
a = 8'd141; b = 8'd17;  #10 
a = 8'd141; b = 8'd18;  #10 
a = 8'd141; b = 8'd19;  #10 
a = 8'd141; b = 8'd20;  #10 
a = 8'd141; b = 8'd21;  #10 
a = 8'd141; b = 8'd22;  #10 
a = 8'd141; b = 8'd23;  #10 
a = 8'd141; b = 8'd24;  #10 
a = 8'd141; b = 8'd25;  #10 
a = 8'd141; b = 8'd26;  #10 
a = 8'd141; b = 8'd27;  #10 
a = 8'd141; b = 8'd28;  #10 
a = 8'd141; b = 8'd29;  #10 
a = 8'd141; b = 8'd30;  #10 
a = 8'd141; b = 8'd31;  #10 
a = 8'd141; b = 8'd32;  #10 
a = 8'd141; b = 8'd33;  #10 
a = 8'd141; b = 8'd34;  #10 
a = 8'd141; b = 8'd35;  #10 
a = 8'd141; b = 8'd36;  #10 
a = 8'd141; b = 8'd37;  #10 
a = 8'd141; b = 8'd38;  #10 
a = 8'd141; b = 8'd39;  #10 
a = 8'd141; b = 8'd40;  #10 
a = 8'd141; b = 8'd41;  #10 
a = 8'd141; b = 8'd42;  #10 
a = 8'd141; b = 8'd43;  #10 
a = 8'd141; b = 8'd44;  #10 
a = 8'd141; b = 8'd45;  #10 
a = 8'd141; b = 8'd46;  #10 
a = 8'd141; b = 8'd47;  #10 
a = 8'd141; b = 8'd48;  #10 
a = 8'd141; b = 8'd49;  #10 
a = 8'd141; b = 8'd50;  #10 
a = 8'd141; b = 8'd51;  #10 
a = 8'd141; b = 8'd52;  #10 
a = 8'd141; b = 8'd53;  #10 
a = 8'd141; b = 8'd54;  #10 
a = 8'd141; b = 8'd55;  #10 
a = 8'd141; b = 8'd56;  #10 
a = 8'd141; b = 8'd57;  #10 
a = 8'd141; b = 8'd58;  #10 
a = 8'd141; b = 8'd59;  #10 
a = 8'd141; b = 8'd60;  #10 
a = 8'd141; b = 8'd61;  #10 
a = 8'd141; b = 8'd62;  #10 
a = 8'd141; b = 8'd63;  #10 
a = 8'd141; b = 8'd64;  #10 
a = 8'd141; b = 8'd65;  #10 
a = 8'd141; b = 8'd66;  #10 
a = 8'd141; b = 8'd67;  #10 
a = 8'd141; b = 8'd68;  #10 
a = 8'd141; b = 8'd69;  #10 
a = 8'd141; b = 8'd70;  #10 
a = 8'd141; b = 8'd71;  #10 
a = 8'd141; b = 8'd72;  #10 
a = 8'd141; b = 8'd73;  #10 
a = 8'd141; b = 8'd74;  #10 
a = 8'd141; b = 8'd75;  #10 
a = 8'd141; b = 8'd76;  #10 
a = 8'd141; b = 8'd77;  #10 
a = 8'd141; b = 8'd78;  #10 
a = 8'd141; b = 8'd79;  #10 
a = 8'd141; b = 8'd80;  #10 
a = 8'd141; b = 8'd81;  #10 
a = 8'd141; b = 8'd82;  #10 
a = 8'd141; b = 8'd83;  #10 
a = 8'd141; b = 8'd84;  #10 
a = 8'd141; b = 8'd85;  #10 
a = 8'd141; b = 8'd86;  #10 
a = 8'd141; b = 8'd87;  #10 
a = 8'd141; b = 8'd88;  #10 
a = 8'd141; b = 8'd89;  #10 
a = 8'd141; b = 8'd90;  #10 
a = 8'd141; b = 8'd91;  #10 
a = 8'd141; b = 8'd92;  #10 
a = 8'd141; b = 8'd93;  #10 
a = 8'd141; b = 8'd94;  #10 
a = 8'd141; b = 8'd95;  #10 
a = 8'd141; b = 8'd96;  #10 
a = 8'd141; b = 8'd97;  #10 
a = 8'd141; b = 8'd98;  #10 
a = 8'd141; b = 8'd99;  #10 
a = 8'd141; b = 8'd100;  #10 
a = 8'd141; b = 8'd101;  #10 
a = 8'd141; b = 8'd102;  #10 
a = 8'd141; b = 8'd103;  #10 
a = 8'd141; b = 8'd104;  #10 
a = 8'd141; b = 8'd105;  #10 
a = 8'd141; b = 8'd106;  #10 
a = 8'd141; b = 8'd107;  #10 
a = 8'd141; b = 8'd108;  #10 
a = 8'd141; b = 8'd109;  #10 
a = 8'd141; b = 8'd110;  #10 
a = 8'd141; b = 8'd111;  #10 
a = 8'd141; b = 8'd112;  #10 
a = 8'd141; b = 8'd113;  #10 
a = 8'd141; b = 8'd114;  #10 
a = 8'd141; b = 8'd115;  #10 
a = 8'd141; b = 8'd116;  #10 
a = 8'd141; b = 8'd117;  #10 
a = 8'd141; b = 8'd118;  #10 
a = 8'd141; b = 8'd119;  #10 
a = 8'd141; b = 8'd120;  #10 
a = 8'd141; b = 8'd121;  #10 
a = 8'd141; b = 8'd122;  #10 
a = 8'd141; b = 8'd123;  #10 
a = 8'd141; b = 8'd124;  #10 
a = 8'd141; b = 8'd125;  #10 
a = 8'd141; b = 8'd126;  #10 
a = 8'd141; b = 8'd127;  #10 
a = 8'd141; b = 8'd128;  #10 
a = 8'd141; b = 8'd129;  #10 
a = 8'd141; b = 8'd130;  #10 
a = 8'd141; b = 8'd131;  #10 
a = 8'd141; b = 8'd132;  #10 
a = 8'd141; b = 8'd133;  #10 
a = 8'd141; b = 8'd134;  #10 
a = 8'd141; b = 8'd135;  #10 
a = 8'd141; b = 8'd136;  #10 
a = 8'd141; b = 8'd137;  #10 
a = 8'd141; b = 8'd138;  #10 
a = 8'd141; b = 8'd139;  #10 
a = 8'd141; b = 8'd140;  #10 
a = 8'd141; b = 8'd141;  #10 
a = 8'd141; b = 8'd142;  #10 
a = 8'd141; b = 8'd143;  #10 
a = 8'd141; b = 8'd144;  #10 
a = 8'd141; b = 8'd145;  #10 
a = 8'd141; b = 8'd146;  #10 
a = 8'd141; b = 8'd147;  #10 
a = 8'd141; b = 8'd148;  #10 
a = 8'd141; b = 8'd149;  #10 
a = 8'd141; b = 8'd150;  #10 
a = 8'd141; b = 8'd151;  #10 
a = 8'd141; b = 8'd152;  #10 
a = 8'd141; b = 8'd153;  #10 
a = 8'd141; b = 8'd154;  #10 
a = 8'd141; b = 8'd155;  #10 
a = 8'd141; b = 8'd156;  #10 
a = 8'd141; b = 8'd157;  #10 
a = 8'd141; b = 8'd158;  #10 
a = 8'd141; b = 8'd159;  #10 
a = 8'd141; b = 8'd160;  #10 
a = 8'd141; b = 8'd161;  #10 
a = 8'd141; b = 8'd162;  #10 
a = 8'd141; b = 8'd163;  #10 
a = 8'd141; b = 8'd164;  #10 
a = 8'd141; b = 8'd165;  #10 
a = 8'd141; b = 8'd166;  #10 
a = 8'd141; b = 8'd167;  #10 
a = 8'd141; b = 8'd168;  #10 
a = 8'd141; b = 8'd169;  #10 
a = 8'd141; b = 8'd170;  #10 
a = 8'd141; b = 8'd171;  #10 
a = 8'd141; b = 8'd172;  #10 
a = 8'd141; b = 8'd173;  #10 
a = 8'd141; b = 8'd174;  #10 
a = 8'd141; b = 8'd175;  #10 
a = 8'd141; b = 8'd176;  #10 
a = 8'd141; b = 8'd177;  #10 
a = 8'd141; b = 8'd178;  #10 
a = 8'd141; b = 8'd179;  #10 
a = 8'd141; b = 8'd180;  #10 
a = 8'd141; b = 8'd181;  #10 
a = 8'd141; b = 8'd182;  #10 
a = 8'd141; b = 8'd183;  #10 
a = 8'd141; b = 8'd184;  #10 
a = 8'd141; b = 8'd185;  #10 
a = 8'd141; b = 8'd186;  #10 
a = 8'd141; b = 8'd187;  #10 
a = 8'd141; b = 8'd188;  #10 
a = 8'd141; b = 8'd189;  #10 
a = 8'd141; b = 8'd190;  #10 
a = 8'd141; b = 8'd191;  #10 
a = 8'd141; b = 8'd192;  #10 
a = 8'd141; b = 8'd193;  #10 
a = 8'd141; b = 8'd194;  #10 
a = 8'd141; b = 8'd195;  #10 
a = 8'd141; b = 8'd196;  #10 
a = 8'd141; b = 8'd197;  #10 
a = 8'd141; b = 8'd198;  #10 
a = 8'd141; b = 8'd199;  #10 
a = 8'd141; b = 8'd200;  #10 
a = 8'd141; b = 8'd201;  #10 
a = 8'd141; b = 8'd202;  #10 
a = 8'd141; b = 8'd203;  #10 
a = 8'd141; b = 8'd204;  #10 
a = 8'd141; b = 8'd205;  #10 
a = 8'd141; b = 8'd206;  #10 
a = 8'd141; b = 8'd207;  #10 
a = 8'd141; b = 8'd208;  #10 
a = 8'd141; b = 8'd209;  #10 
a = 8'd141; b = 8'd210;  #10 
a = 8'd141; b = 8'd211;  #10 
a = 8'd141; b = 8'd212;  #10 
a = 8'd141; b = 8'd213;  #10 
a = 8'd141; b = 8'd214;  #10 
a = 8'd141; b = 8'd215;  #10 
a = 8'd141; b = 8'd216;  #10 
a = 8'd141; b = 8'd217;  #10 
a = 8'd141; b = 8'd218;  #10 
a = 8'd141; b = 8'd219;  #10 
a = 8'd141; b = 8'd220;  #10 
a = 8'd141; b = 8'd221;  #10 
a = 8'd141; b = 8'd222;  #10 
a = 8'd141; b = 8'd223;  #10 
a = 8'd141; b = 8'd224;  #10 
a = 8'd141; b = 8'd225;  #10 
a = 8'd141; b = 8'd226;  #10 
a = 8'd141; b = 8'd227;  #10 
a = 8'd141; b = 8'd228;  #10 
a = 8'd141; b = 8'd229;  #10 
a = 8'd141; b = 8'd230;  #10 
a = 8'd141; b = 8'd231;  #10 
a = 8'd141; b = 8'd232;  #10 
a = 8'd141; b = 8'd233;  #10 
a = 8'd141; b = 8'd234;  #10 
a = 8'd141; b = 8'd235;  #10 
a = 8'd141; b = 8'd236;  #10 
a = 8'd141; b = 8'd237;  #10 
a = 8'd141; b = 8'd238;  #10 
a = 8'd141; b = 8'd239;  #10 
a = 8'd141; b = 8'd240;  #10 
a = 8'd141; b = 8'd241;  #10 
a = 8'd141; b = 8'd242;  #10 
a = 8'd141; b = 8'd243;  #10 
a = 8'd141; b = 8'd244;  #10 
a = 8'd141; b = 8'd245;  #10 
a = 8'd141; b = 8'd246;  #10 
a = 8'd141; b = 8'd247;  #10 
a = 8'd141; b = 8'd248;  #10 
a = 8'd141; b = 8'd249;  #10 
a = 8'd141; b = 8'd250;  #10 
a = 8'd141; b = 8'd251;  #10 
a = 8'd141; b = 8'd252;  #10 
a = 8'd141; b = 8'd253;  #10 
a = 8'd141; b = 8'd254;  #10 
a = 8'd141; b = 8'd255;  #10 
a = 8'd142; b = 8'd0;  #10 
a = 8'd142; b = 8'd1;  #10 
a = 8'd142; b = 8'd2;  #10 
a = 8'd142; b = 8'd3;  #10 
a = 8'd142; b = 8'd4;  #10 
a = 8'd142; b = 8'd5;  #10 
a = 8'd142; b = 8'd6;  #10 
a = 8'd142; b = 8'd7;  #10 
a = 8'd142; b = 8'd8;  #10 
a = 8'd142; b = 8'd9;  #10 
a = 8'd142; b = 8'd10;  #10 
a = 8'd142; b = 8'd11;  #10 
a = 8'd142; b = 8'd12;  #10 
a = 8'd142; b = 8'd13;  #10 
a = 8'd142; b = 8'd14;  #10 
a = 8'd142; b = 8'd15;  #10 
a = 8'd142; b = 8'd16;  #10 
a = 8'd142; b = 8'd17;  #10 
a = 8'd142; b = 8'd18;  #10 
a = 8'd142; b = 8'd19;  #10 
a = 8'd142; b = 8'd20;  #10 
a = 8'd142; b = 8'd21;  #10 
a = 8'd142; b = 8'd22;  #10 
a = 8'd142; b = 8'd23;  #10 
a = 8'd142; b = 8'd24;  #10 
a = 8'd142; b = 8'd25;  #10 
a = 8'd142; b = 8'd26;  #10 
a = 8'd142; b = 8'd27;  #10 
a = 8'd142; b = 8'd28;  #10 
a = 8'd142; b = 8'd29;  #10 
a = 8'd142; b = 8'd30;  #10 
a = 8'd142; b = 8'd31;  #10 
a = 8'd142; b = 8'd32;  #10 
a = 8'd142; b = 8'd33;  #10 
a = 8'd142; b = 8'd34;  #10 
a = 8'd142; b = 8'd35;  #10 
a = 8'd142; b = 8'd36;  #10 
a = 8'd142; b = 8'd37;  #10 
a = 8'd142; b = 8'd38;  #10 
a = 8'd142; b = 8'd39;  #10 
a = 8'd142; b = 8'd40;  #10 
a = 8'd142; b = 8'd41;  #10 
a = 8'd142; b = 8'd42;  #10 
a = 8'd142; b = 8'd43;  #10 
a = 8'd142; b = 8'd44;  #10 
a = 8'd142; b = 8'd45;  #10 
a = 8'd142; b = 8'd46;  #10 
a = 8'd142; b = 8'd47;  #10 
a = 8'd142; b = 8'd48;  #10 
a = 8'd142; b = 8'd49;  #10 
a = 8'd142; b = 8'd50;  #10 
a = 8'd142; b = 8'd51;  #10 
a = 8'd142; b = 8'd52;  #10 
a = 8'd142; b = 8'd53;  #10 
a = 8'd142; b = 8'd54;  #10 
a = 8'd142; b = 8'd55;  #10 
a = 8'd142; b = 8'd56;  #10 
a = 8'd142; b = 8'd57;  #10 
a = 8'd142; b = 8'd58;  #10 
a = 8'd142; b = 8'd59;  #10 
a = 8'd142; b = 8'd60;  #10 
a = 8'd142; b = 8'd61;  #10 
a = 8'd142; b = 8'd62;  #10 
a = 8'd142; b = 8'd63;  #10 
a = 8'd142; b = 8'd64;  #10 
a = 8'd142; b = 8'd65;  #10 
a = 8'd142; b = 8'd66;  #10 
a = 8'd142; b = 8'd67;  #10 
a = 8'd142; b = 8'd68;  #10 
a = 8'd142; b = 8'd69;  #10 
a = 8'd142; b = 8'd70;  #10 
a = 8'd142; b = 8'd71;  #10 
a = 8'd142; b = 8'd72;  #10 
a = 8'd142; b = 8'd73;  #10 
a = 8'd142; b = 8'd74;  #10 
a = 8'd142; b = 8'd75;  #10 
a = 8'd142; b = 8'd76;  #10 
a = 8'd142; b = 8'd77;  #10 
a = 8'd142; b = 8'd78;  #10 
a = 8'd142; b = 8'd79;  #10 
a = 8'd142; b = 8'd80;  #10 
a = 8'd142; b = 8'd81;  #10 
a = 8'd142; b = 8'd82;  #10 
a = 8'd142; b = 8'd83;  #10 
a = 8'd142; b = 8'd84;  #10 
a = 8'd142; b = 8'd85;  #10 
a = 8'd142; b = 8'd86;  #10 
a = 8'd142; b = 8'd87;  #10 
a = 8'd142; b = 8'd88;  #10 
a = 8'd142; b = 8'd89;  #10 
a = 8'd142; b = 8'd90;  #10 
a = 8'd142; b = 8'd91;  #10 
a = 8'd142; b = 8'd92;  #10 
a = 8'd142; b = 8'd93;  #10 
a = 8'd142; b = 8'd94;  #10 
a = 8'd142; b = 8'd95;  #10 
a = 8'd142; b = 8'd96;  #10 
a = 8'd142; b = 8'd97;  #10 
a = 8'd142; b = 8'd98;  #10 
a = 8'd142; b = 8'd99;  #10 
a = 8'd142; b = 8'd100;  #10 
a = 8'd142; b = 8'd101;  #10 
a = 8'd142; b = 8'd102;  #10 
a = 8'd142; b = 8'd103;  #10 
a = 8'd142; b = 8'd104;  #10 
a = 8'd142; b = 8'd105;  #10 
a = 8'd142; b = 8'd106;  #10 
a = 8'd142; b = 8'd107;  #10 
a = 8'd142; b = 8'd108;  #10 
a = 8'd142; b = 8'd109;  #10 
a = 8'd142; b = 8'd110;  #10 
a = 8'd142; b = 8'd111;  #10 
a = 8'd142; b = 8'd112;  #10 
a = 8'd142; b = 8'd113;  #10 
a = 8'd142; b = 8'd114;  #10 
a = 8'd142; b = 8'd115;  #10 
a = 8'd142; b = 8'd116;  #10 
a = 8'd142; b = 8'd117;  #10 
a = 8'd142; b = 8'd118;  #10 
a = 8'd142; b = 8'd119;  #10 
a = 8'd142; b = 8'd120;  #10 
a = 8'd142; b = 8'd121;  #10 
a = 8'd142; b = 8'd122;  #10 
a = 8'd142; b = 8'd123;  #10 
a = 8'd142; b = 8'd124;  #10 
a = 8'd142; b = 8'd125;  #10 
a = 8'd142; b = 8'd126;  #10 
a = 8'd142; b = 8'd127;  #10 
a = 8'd142; b = 8'd128;  #10 
a = 8'd142; b = 8'd129;  #10 
a = 8'd142; b = 8'd130;  #10 
a = 8'd142; b = 8'd131;  #10 
a = 8'd142; b = 8'd132;  #10 
a = 8'd142; b = 8'd133;  #10 
a = 8'd142; b = 8'd134;  #10 
a = 8'd142; b = 8'd135;  #10 
a = 8'd142; b = 8'd136;  #10 
a = 8'd142; b = 8'd137;  #10 
a = 8'd142; b = 8'd138;  #10 
a = 8'd142; b = 8'd139;  #10 
a = 8'd142; b = 8'd140;  #10 
a = 8'd142; b = 8'd141;  #10 
a = 8'd142; b = 8'd142;  #10 
a = 8'd142; b = 8'd143;  #10 
a = 8'd142; b = 8'd144;  #10 
a = 8'd142; b = 8'd145;  #10 
a = 8'd142; b = 8'd146;  #10 
a = 8'd142; b = 8'd147;  #10 
a = 8'd142; b = 8'd148;  #10 
a = 8'd142; b = 8'd149;  #10 
a = 8'd142; b = 8'd150;  #10 
a = 8'd142; b = 8'd151;  #10 
a = 8'd142; b = 8'd152;  #10 
a = 8'd142; b = 8'd153;  #10 
a = 8'd142; b = 8'd154;  #10 
a = 8'd142; b = 8'd155;  #10 
a = 8'd142; b = 8'd156;  #10 
a = 8'd142; b = 8'd157;  #10 
a = 8'd142; b = 8'd158;  #10 
a = 8'd142; b = 8'd159;  #10 
a = 8'd142; b = 8'd160;  #10 
a = 8'd142; b = 8'd161;  #10 
a = 8'd142; b = 8'd162;  #10 
a = 8'd142; b = 8'd163;  #10 
a = 8'd142; b = 8'd164;  #10 
a = 8'd142; b = 8'd165;  #10 
a = 8'd142; b = 8'd166;  #10 
a = 8'd142; b = 8'd167;  #10 
a = 8'd142; b = 8'd168;  #10 
a = 8'd142; b = 8'd169;  #10 
a = 8'd142; b = 8'd170;  #10 
a = 8'd142; b = 8'd171;  #10 
a = 8'd142; b = 8'd172;  #10 
a = 8'd142; b = 8'd173;  #10 
a = 8'd142; b = 8'd174;  #10 
a = 8'd142; b = 8'd175;  #10 
a = 8'd142; b = 8'd176;  #10 
a = 8'd142; b = 8'd177;  #10 
a = 8'd142; b = 8'd178;  #10 
a = 8'd142; b = 8'd179;  #10 
a = 8'd142; b = 8'd180;  #10 
a = 8'd142; b = 8'd181;  #10 
a = 8'd142; b = 8'd182;  #10 
a = 8'd142; b = 8'd183;  #10 
a = 8'd142; b = 8'd184;  #10 
a = 8'd142; b = 8'd185;  #10 
a = 8'd142; b = 8'd186;  #10 
a = 8'd142; b = 8'd187;  #10 
a = 8'd142; b = 8'd188;  #10 
a = 8'd142; b = 8'd189;  #10 
a = 8'd142; b = 8'd190;  #10 
a = 8'd142; b = 8'd191;  #10 
a = 8'd142; b = 8'd192;  #10 
a = 8'd142; b = 8'd193;  #10 
a = 8'd142; b = 8'd194;  #10 
a = 8'd142; b = 8'd195;  #10 
a = 8'd142; b = 8'd196;  #10 
a = 8'd142; b = 8'd197;  #10 
a = 8'd142; b = 8'd198;  #10 
a = 8'd142; b = 8'd199;  #10 
a = 8'd142; b = 8'd200;  #10 
a = 8'd142; b = 8'd201;  #10 
a = 8'd142; b = 8'd202;  #10 
a = 8'd142; b = 8'd203;  #10 
a = 8'd142; b = 8'd204;  #10 
a = 8'd142; b = 8'd205;  #10 
a = 8'd142; b = 8'd206;  #10 
a = 8'd142; b = 8'd207;  #10 
a = 8'd142; b = 8'd208;  #10 
a = 8'd142; b = 8'd209;  #10 
a = 8'd142; b = 8'd210;  #10 
a = 8'd142; b = 8'd211;  #10 
a = 8'd142; b = 8'd212;  #10 
a = 8'd142; b = 8'd213;  #10 
a = 8'd142; b = 8'd214;  #10 
a = 8'd142; b = 8'd215;  #10 
a = 8'd142; b = 8'd216;  #10 
a = 8'd142; b = 8'd217;  #10 
a = 8'd142; b = 8'd218;  #10 
a = 8'd142; b = 8'd219;  #10 
a = 8'd142; b = 8'd220;  #10 
a = 8'd142; b = 8'd221;  #10 
a = 8'd142; b = 8'd222;  #10 
a = 8'd142; b = 8'd223;  #10 
a = 8'd142; b = 8'd224;  #10 
a = 8'd142; b = 8'd225;  #10 
a = 8'd142; b = 8'd226;  #10 
a = 8'd142; b = 8'd227;  #10 
a = 8'd142; b = 8'd228;  #10 
a = 8'd142; b = 8'd229;  #10 
a = 8'd142; b = 8'd230;  #10 
a = 8'd142; b = 8'd231;  #10 
a = 8'd142; b = 8'd232;  #10 
a = 8'd142; b = 8'd233;  #10 
a = 8'd142; b = 8'd234;  #10 
a = 8'd142; b = 8'd235;  #10 
a = 8'd142; b = 8'd236;  #10 
a = 8'd142; b = 8'd237;  #10 
a = 8'd142; b = 8'd238;  #10 
a = 8'd142; b = 8'd239;  #10 
a = 8'd142; b = 8'd240;  #10 
a = 8'd142; b = 8'd241;  #10 
a = 8'd142; b = 8'd242;  #10 
a = 8'd142; b = 8'd243;  #10 
a = 8'd142; b = 8'd244;  #10 
a = 8'd142; b = 8'd245;  #10 
a = 8'd142; b = 8'd246;  #10 
a = 8'd142; b = 8'd247;  #10 
a = 8'd142; b = 8'd248;  #10 
a = 8'd142; b = 8'd249;  #10 
a = 8'd142; b = 8'd250;  #10 
a = 8'd142; b = 8'd251;  #10 
a = 8'd142; b = 8'd252;  #10 
a = 8'd142; b = 8'd253;  #10 
a = 8'd142; b = 8'd254;  #10 
a = 8'd142; b = 8'd255;  #10 
a = 8'd143; b = 8'd0;  #10 
a = 8'd143; b = 8'd1;  #10 
a = 8'd143; b = 8'd2;  #10 
a = 8'd143; b = 8'd3;  #10 
a = 8'd143; b = 8'd4;  #10 
a = 8'd143; b = 8'd5;  #10 
a = 8'd143; b = 8'd6;  #10 
a = 8'd143; b = 8'd7;  #10 
a = 8'd143; b = 8'd8;  #10 
a = 8'd143; b = 8'd9;  #10 
a = 8'd143; b = 8'd10;  #10 
a = 8'd143; b = 8'd11;  #10 
a = 8'd143; b = 8'd12;  #10 
a = 8'd143; b = 8'd13;  #10 
a = 8'd143; b = 8'd14;  #10 
a = 8'd143; b = 8'd15;  #10 
a = 8'd143; b = 8'd16;  #10 
a = 8'd143; b = 8'd17;  #10 
a = 8'd143; b = 8'd18;  #10 
a = 8'd143; b = 8'd19;  #10 
a = 8'd143; b = 8'd20;  #10 
a = 8'd143; b = 8'd21;  #10 
a = 8'd143; b = 8'd22;  #10 
a = 8'd143; b = 8'd23;  #10 
a = 8'd143; b = 8'd24;  #10 
a = 8'd143; b = 8'd25;  #10 
a = 8'd143; b = 8'd26;  #10 
a = 8'd143; b = 8'd27;  #10 
a = 8'd143; b = 8'd28;  #10 
a = 8'd143; b = 8'd29;  #10 
a = 8'd143; b = 8'd30;  #10 
a = 8'd143; b = 8'd31;  #10 
a = 8'd143; b = 8'd32;  #10 
a = 8'd143; b = 8'd33;  #10 
a = 8'd143; b = 8'd34;  #10 
a = 8'd143; b = 8'd35;  #10 
a = 8'd143; b = 8'd36;  #10 
a = 8'd143; b = 8'd37;  #10 
a = 8'd143; b = 8'd38;  #10 
a = 8'd143; b = 8'd39;  #10 
a = 8'd143; b = 8'd40;  #10 
a = 8'd143; b = 8'd41;  #10 
a = 8'd143; b = 8'd42;  #10 
a = 8'd143; b = 8'd43;  #10 
a = 8'd143; b = 8'd44;  #10 
a = 8'd143; b = 8'd45;  #10 
a = 8'd143; b = 8'd46;  #10 
a = 8'd143; b = 8'd47;  #10 
a = 8'd143; b = 8'd48;  #10 
a = 8'd143; b = 8'd49;  #10 
a = 8'd143; b = 8'd50;  #10 
a = 8'd143; b = 8'd51;  #10 
a = 8'd143; b = 8'd52;  #10 
a = 8'd143; b = 8'd53;  #10 
a = 8'd143; b = 8'd54;  #10 
a = 8'd143; b = 8'd55;  #10 
a = 8'd143; b = 8'd56;  #10 
a = 8'd143; b = 8'd57;  #10 
a = 8'd143; b = 8'd58;  #10 
a = 8'd143; b = 8'd59;  #10 
a = 8'd143; b = 8'd60;  #10 
a = 8'd143; b = 8'd61;  #10 
a = 8'd143; b = 8'd62;  #10 
a = 8'd143; b = 8'd63;  #10 
a = 8'd143; b = 8'd64;  #10 
a = 8'd143; b = 8'd65;  #10 
a = 8'd143; b = 8'd66;  #10 
a = 8'd143; b = 8'd67;  #10 
a = 8'd143; b = 8'd68;  #10 
a = 8'd143; b = 8'd69;  #10 
a = 8'd143; b = 8'd70;  #10 
a = 8'd143; b = 8'd71;  #10 
a = 8'd143; b = 8'd72;  #10 
a = 8'd143; b = 8'd73;  #10 
a = 8'd143; b = 8'd74;  #10 
a = 8'd143; b = 8'd75;  #10 
a = 8'd143; b = 8'd76;  #10 
a = 8'd143; b = 8'd77;  #10 
a = 8'd143; b = 8'd78;  #10 
a = 8'd143; b = 8'd79;  #10 
a = 8'd143; b = 8'd80;  #10 
a = 8'd143; b = 8'd81;  #10 
a = 8'd143; b = 8'd82;  #10 
a = 8'd143; b = 8'd83;  #10 
a = 8'd143; b = 8'd84;  #10 
a = 8'd143; b = 8'd85;  #10 
a = 8'd143; b = 8'd86;  #10 
a = 8'd143; b = 8'd87;  #10 
a = 8'd143; b = 8'd88;  #10 
a = 8'd143; b = 8'd89;  #10 
a = 8'd143; b = 8'd90;  #10 
a = 8'd143; b = 8'd91;  #10 
a = 8'd143; b = 8'd92;  #10 
a = 8'd143; b = 8'd93;  #10 
a = 8'd143; b = 8'd94;  #10 
a = 8'd143; b = 8'd95;  #10 
a = 8'd143; b = 8'd96;  #10 
a = 8'd143; b = 8'd97;  #10 
a = 8'd143; b = 8'd98;  #10 
a = 8'd143; b = 8'd99;  #10 
a = 8'd143; b = 8'd100;  #10 
a = 8'd143; b = 8'd101;  #10 
a = 8'd143; b = 8'd102;  #10 
a = 8'd143; b = 8'd103;  #10 
a = 8'd143; b = 8'd104;  #10 
a = 8'd143; b = 8'd105;  #10 
a = 8'd143; b = 8'd106;  #10 
a = 8'd143; b = 8'd107;  #10 
a = 8'd143; b = 8'd108;  #10 
a = 8'd143; b = 8'd109;  #10 
a = 8'd143; b = 8'd110;  #10 
a = 8'd143; b = 8'd111;  #10 
a = 8'd143; b = 8'd112;  #10 
a = 8'd143; b = 8'd113;  #10 
a = 8'd143; b = 8'd114;  #10 
a = 8'd143; b = 8'd115;  #10 
a = 8'd143; b = 8'd116;  #10 
a = 8'd143; b = 8'd117;  #10 
a = 8'd143; b = 8'd118;  #10 
a = 8'd143; b = 8'd119;  #10 
a = 8'd143; b = 8'd120;  #10 
a = 8'd143; b = 8'd121;  #10 
a = 8'd143; b = 8'd122;  #10 
a = 8'd143; b = 8'd123;  #10 
a = 8'd143; b = 8'd124;  #10 
a = 8'd143; b = 8'd125;  #10 
a = 8'd143; b = 8'd126;  #10 
a = 8'd143; b = 8'd127;  #10 
a = 8'd143; b = 8'd128;  #10 
a = 8'd143; b = 8'd129;  #10 
a = 8'd143; b = 8'd130;  #10 
a = 8'd143; b = 8'd131;  #10 
a = 8'd143; b = 8'd132;  #10 
a = 8'd143; b = 8'd133;  #10 
a = 8'd143; b = 8'd134;  #10 
a = 8'd143; b = 8'd135;  #10 
a = 8'd143; b = 8'd136;  #10 
a = 8'd143; b = 8'd137;  #10 
a = 8'd143; b = 8'd138;  #10 
a = 8'd143; b = 8'd139;  #10 
a = 8'd143; b = 8'd140;  #10 
a = 8'd143; b = 8'd141;  #10 
a = 8'd143; b = 8'd142;  #10 
a = 8'd143; b = 8'd143;  #10 
a = 8'd143; b = 8'd144;  #10 
a = 8'd143; b = 8'd145;  #10 
a = 8'd143; b = 8'd146;  #10 
a = 8'd143; b = 8'd147;  #10 
a = 8'd143; b = 8'd148;  #10 
a = 8'd143; b = 8'd149;  #10 
a = 8'd143; b = 8'd150;  #10 
a = 8'd143; b = 8'd151;  #10 
a = 8'd143; b = 8'd152;  #10 
a = 8'd143; b = 8'd153;  #10 
a = 8'd143; b = 8'd154;  #10 
a = 8'd143; b = 8'd155;  #10 
a = 8'd143; b = 8'd156;  #10 
a = 8'd143; b = 8'd157;  #10 
a = 8'd143; b = 8'd158;  #10 
a = 8'd143; b = 8'd159;  #10 
a = 8'd143; b = 8'd160;  #10 
a = 8'd143; b = 8'd161;  #10 
a = 8'd143; b = 8'd162;  #10 
a = 8'd143; b = 8'd163;  #10 
a = 8'd143; b = 8'd164;  #10 
a = 8'd143; b = 8'd165;  #10 
a = 8'd143; b = 8'd166;  #10 
a = 8'd143; b = 8'd167;  #10 
a = 8'd143; b = 8'd168;  #10 
a = 8'd143; b = 8'd169;  #10 
a = 8'd143; b = 8'd170;  #10 
a = 8'd143; b = 8'd171;  #10 
a = 8'd143; b = 8'd172;  #10 
a = 8'd143; b = 8'd173;  #10 
a = 8'd143; b = 8'd174;  #10 
a = 8'd143; b = 8'd175;  #10 
a = 8'd143; b = 8'd176;  #10 
a = 8'd143; b = 8'd177;  #10 
a = 8'd143; b = 8'd178;  #10 
a = 8'd143; b = 8'd179;  #10 
a = 8'd143; b = 8'd180;  #10 
a = 8'd143; b = 8'd181;  #10 
a = 8'd143; b = 8'd182;  #10 
a = 8'd143; b = 8'd183;  #10 
a = 8'd143; b = 8'd184;  #10 
a = 8'd143; b = 8'd185;  #10 
a = 8'd143; b = 8'd186;  #10 
a = 8'd143; b = 8'd187;  #10 
a = 8'd143; b = 8'd188;  #10 
a = 8'd143; b = 8'd189;  #10 
a = 8'd143; b = 8'd190;  #10 
a = 8'd143; b = 8'd191;  #10 
a = 8'd143; b = 8'd192;  #10 
a = 8'd143; b = 8'd193;  #10 
a = 8'd143; b = 8'd194;  #10 
a = 8'd143; b = 8'd195;  #10 
a = 8'd143; b = 8'd196;  #10 
a = 8'd143; b = 8'd197;  #10 
a = 8'd143; b = 8'd198;  #10 
a = 8'd143; b = 8'd199;  #10 
a = 8'd143; b = 8'd200;  #10 
a = 8'd143; b = 8'd201;  #10 
a = 8'd143; b = 8'd202;  #10 
a = 8'd143; b = 8'd203;  #10 
a = 8'd143; b = 8'd204;  #10 
a = 8'd143; b = 8'd205;  #10 
a = 8'd143; b = 8'd206;  #10 
a = 8'd143; b = 8'd207;  #10 
a = 8'd143; b = 8'd208;  #10 
a = 8'd143; b = 8'd209;  #10 
a = 8'd143; b = 8'd210;  #10 
a = 8'd143; b = 8'd211;  #10 
a = 8'd143; b = 8'd212;  #10 
a = 8'd143; b = 8'd213;  #10 
a = 8'd143; b = 8'd214;  #10 
a = 8'd143; b = 8'd215;  #10 
a = 8'd143; b = 8'd216;  #10 
a = 8'd143; b = 8'd217;  #10 
a = 8'd143; b = 8'd218;  #10 
a = 8'd143; b = 8'd219;  #10 
a = 8'd143; b = 8'd220;  #10 
a = 8'd143; b = 8'd221;  #10 
a = 8'd143; b = 8'd222;  #10 
a = 8'd143; b = 8'd223;  #10 
a = 8'd143; b = 8'd224;  #10 
a = 8'd143; b = 8'd225;  #10 
a = 8'd143; b = 8'd226;  #10 
a = 8'd143; b = 8'd227;  #10 
a = 8'd143; b = 8'd228;  #10 
a = 8'd143; b = 8'd229;  #10 
a = 8'd143; b = 8'd230;  #10 
a = 8'd143; b = 8'd231;  #10 
a = 8'd143; b = 8'd232;  #10 
a = 8'd143; b = 8'd233;  #10 
a = 8'd143; b = 8'd234;  #10 
a = 8'd143; b = 8'd235;  #10 
a = 8'd143; b = 8'd236;  #10 
a = 8'd143; b = 8'd237;  #10 
a = 8'd143; b = 8'd238;  #10 
a = 8'd143; b = 8'd239;  #10 
a = 8'd143; b = 8'd240;  #10 
a = 8'd143; b = 8'd241;  #10 
a = 8'd143; b = 8'd242;  #10 
a = 8'd143; b = 8'd243;  #10 
a = 8'd143; b = 8'd244;  #10 
a = 8'd143; b = 8'd245;  #10 
a = 8'd143; b = 8'd246;  #10 
a = 8'd143; b = 8'd247;  #10 
a = 8'd143; b = 8'd248;  #10 
a = 8'd143; b = 8'd249;  #10 
a = 8'd143; b = 8'd250;  #10 
a = 8'd143; b = 8'd251;  #10 
a = 8'd143; b = 8'd252;  #10 
a = 8'd143; b = 8'd253;  #10 
a = 8'd143; b = 8'd254;  #10 
a = 8'd143; b = 8'd255;  #10 
a = 8'd144; b = 8'd0;  #10 
a = 8'd144; b = 8'd1;  #10 
a = 8'd144; b = 8'd2;  #10 
a = 8'd144; b = 8'd3;  #10 
a = 8'd144; b = 8'd4;  #10 
a = 8'd144; b = 8'd5;  #10 
a = 8'd144; b = 8'd6;  #10 
a = 8'd144; b = 8'd7;  #10 
a = 8'd144; b = 8'd8;  #10 
a = 8'd144; b = 8'd9;  #10 
a = 8'd144; b = 8'd10;  #10 
a = 8'd144; b = 8'd11;  #10 
a = 8'd144; b = 8'd12;  #10 
a = 8'd144; b = 8'd13;  #10 
a = 8'd144; b = 8'd14;  #10 
a = 8'd144; b = 8'd15;  #10 
a = 8'd144; b = 8'd16;  #10 
a = 8'd144; b = 8'd17;  #10 
a = 8'd144; b = 8'd18;  #10 
a = 8'd144; b = 8'd19;  #10 
a = 8'd144; b = 8'd20;  #10 
a = 8'd144; b = 8'd21;  #10 
a = 8'd144; b = 8'd22;  #10 
a = 8'd144; b = 8'd23;  #10 
a = 8'd144; b = 8'd24;  #10 
a = 8'd144; b = 8'd25;  #10 
a = 8'd144; b = 8'd26;  #10 
a = 8'd144; b = 8'd27;  #10 
a = 8'd144; b = 8'd28;  #10 
a = 8'd144; b = 8'd29;  #10 
a = 8'd144; b = 8'd30;  #10 
a = 8'd144; b = 8'd31;  #10 
a = 8'd144; b = 8'd32;  #10 
a = 8'd144; b = 8'd33;  #10 
a = 8'd144; b = 8'd34;  #10 
a = 8'd144; b = 8'd35;  #10 
a = 8'd144; b = 8'd36;  #10 
a = 8'd144; b = 8'd37;  #10 
a = 8'd144; b = 8'd38;  #10 
a = 8'd144; b = 8'd39;  #10 
a = 8'd144; b = 8'd40;  #10 
a = 8'd144; b = 8'd41;  #10 
a = 8'd144; b = 8'd42;  #10 
a = 8'd144; b = 8'd43;  #10 
a = 8'd144; b = 8'd44;  #10 
a = 8'd144; b = 8'd45;  #10 
a = 8'd144; b = 8'd46;  #10 
a = 8'd144; b = 8'd47;  #10 
a = 8'd144; b = 8'd48;  #10 
a = 8'd144; b = 8'd49;  #10 
a = 8'd144; b = 8'd50;  #10 
a = 8'd144; b = 8'd51;  #10 
a = 8'd144; b = 8'd52;  #10 
a = 8'd144; b = 8'd53;  #10 
a = 8'd144; b = 8'd54;  #10 
a = 8'd144; b = 8'd55;  #10 
a = 8'd144; b = 8'd56;  #10 
a = 8'd144; b = 8'd57;  #10 
a = 8'd144; b = 8'd58;  #10 
a = 8'd144; b = 8'd59;  #10 
a = 8'd144; b = 8'd60;  #10 
a = 8'd144; b = 8'd61;  #10 
a = 8'd144; b = 8'd62;  #10 
a = 8'd144; b = 8'd63;  #10 
a = 8'd144; b = 8'd64;  #10 
a = 8'd144; b = 8'd65;  #10 
a = 8'd144; b = 8'd66;  #10 
a = 8'd144; b = 8'd67;  #10 
a = 8'd144; b = 8'd68;  #10 
a = 8'd144; b = 8'd69;  #10 
a = 8'd144; b = 8'd70;  #10 
a = 8'd144; b = 8'd71;  #10 
a = 8'd144; b = 8'd72;  #10 
a = 8'd144; b = 8'd73;  #10 
a = 8'd144; b = 8'd74;  #10 
a = 8'd144; b = 8'd75;  #10 
a = 8'd144; b = 8'd76;  #10 
a = 8'd144; b = 8'd77;  #10 
a = 8'd144; b = 8'd78;  #10 
a = 8'd144; b = 8'd79;  #10 
a = 8'd144; b = 8'd80;  #10 
a = 8'd144; b = 8'd81;  #10 
a = 8'd144; b = 8'd82;  #10 
a = 8'd144; b = 8'd83;  #10 
a = 8'd144; b = 8'd84;  #10 
a = 8'd144; b = 8'd85;  #10 
a = 8'd144; b = 8'd86;  #10 
a = 8'd144; b = 8'd87;  #10 
a = 8'd144; b = 8'd88;  #10 
a = 8'd144; b = 8'd89;  #10 
a = 8'd144; b = 8'd90;  #10 
a = 8'd144; b = 8'd91;  #10 
a = 8'd144; b = 8'd92;  #10 
a = 8'd144; b = 8'd93;  #10 
a = 8'd144; b = 8'd94;  #10 
a = 8'd144; b = 8'd95;  #10 
a = 8'd144; b = 8'd96;  #10 
a = 8'd144; b = 8'd97;  #10 
a = 8'd144; b = 8'd98;  #10 
a = 8'd144; b = 8'd99;  #10 
a = 8'd144; b = 8'd100;  #10 
a = 8'd144; b = 8'd101;  #10 
a = 8'd144; b = 8'd102;  #10 
a = 8'd144; b = 8'd103;  #10 
a = 8'd144; b = 8'd104;  #10 
a = 8'd144; b = 8'd105;  #10 
a = 8'd144; b = 8'd106;  #10 
a = 8'd144; b = 8'd107;  #10 
a = 8'd144; b = 8'd108;  #10 
a = 8'd144; b = 8'd109;  #10 
a = 8'd144; b = 8'd110;  #10 
a = 8'd144; b = 8'd111;  #10 
a = 8'd144; b = 8'd112;  #10 
a = 8'd144; b = 8'd113;  #10 
a = 8'd144; b = 8'd114;  #10 
a = 8'd144; b = 8'd115;  #10 
a = 8'd144; b = 8'd116;  #10 
a = 8'd144; b = 8'd117;  #10 
a = 8'd144; b = 8'd118;  #10 
a = 8'd144; b = 8'd119;  #10 
a = 8'd144; b = 8'd120;  #10 
a = 8'd144; b = 8'd121;  #10 
a = 8'd144; b = 8'd122;  #10 
a = 8'd144; b = 8'd123;  #10 
a = 8'd144; b = 8'd124;  #10 
a = 8'd144; b = 8'd125;  #10 
a = 8'd144; b = 8'd126;  #10 
a = 8'd144; b = 8'd127;  #10 
a = 8'd144; b = 8'd128;  #10 
a = 8'd144; b = 8'd129;  #10 
a = 8'd144; b = 8'd130;  #10 
a = 8'd144; b = 8'd131;  #10 
a = 8'd144; b = 8'd132;  #10 
a = 8'd144; b = 8'd133;  #10 
a = 8'd144; b = 8'd134;  #10 
a = 8'd144; b = 8'd135;  #10 
a = 8'd144; b = 8'd136;  #10 
a = 8'd144; b = 8'd137;  #10 
a = 8'd144; b = 8'd138;  #10 
a = 8'd144; b = 8'd139;  #10 
a = 8'd144; b = 8'd140;  #10 
a = 8'd144; b = 8'd141;  #10 
a = 8'd144; b = 8'd142;  #10 
a = 8'd144; b = 8'd143;  #10 
a = 8'd144; b = 8'd144;  #10 
a = 8'd144; b = 8'd145;  #10 
a = 8'd144; b = 8'd146;  #10 
a = 8'd144; b = 8'd147;  #10 
a = 8'd144; b = 8'd148;  #10 
a = 8'd144; b = 8'd149;  #10 
a = 8'd144; b = 8'd150;  #10 
a = 8'd144; b = 8'd151;  #10 
a = 8'd144; b = 8'd152;  #10 
a = 8'd144; b = 8'd153;  #10 
a = 8'd144; b = 8'd154;  #10 
a = 8'd144; b = 8'd155;  #10 
a = 8'd144; b = 8'd156;  #10 
a = 8'd144; b = 8'd157;  #10 
a = 8'd144; b = 8'd158;  #10 
a = 8'd144; b = 8'd159;  #10 
a = 8'd144; b = 8'd160;  #10 
a = 8'd144; b = 8'd161;  #10 
a = 8'd144; b = 8'd162;  #10 
a = 8'd144; b = 8'd163;  #10 
a = 8'd144; b = 8'd164;  #10 
a = 8'd144; b = 8'd165;  #10 
a = 8'd144; b = 8'd166;  #10 
a = 8'd144; b = 8'd167;  #10 
a = 8'd144; b = 8'd168;  #10 
a = 8'd144; b = 8'd169;  #10 
a = 8'd144; b = 8'd170;  #10 
a = 8'd144; b = 8'd171;  #10 
a = 8'd144; b = 8'd172;  #10 
a = 8'd144; b = 8'd173;  #10 
a = 8'd144; b = 8'd174;  #10 
a = 8'd144; b = 8'd175;  #10 
a = 8'd144; b = 8'd176;  #10 
a = 8'd144; b = 8'd177;  #10 
a = 8'd144; b = 8'd178;  #10 
a = 8'd144; b = 8'd179;  #10 
a = 8'd144; b = 8'd180;  #10 
a = 8'd144; b = 8'd181;  #10 
a = 8'd144; b = 8'd182;  #10 
a = 8'd144; b = 8'd183;  #10 
a = 8'd144; b = 8'd184;  #10 
a = 8'd144; b = 8'd185;  #10 
a = 8'd144; b = 8'd186;  #10 
a = 8'd144; b = 8'd187;  #10 
a = 8'd144; b = 8'd188;  #10 
a = 8'd144; b = 8'd189;  #10 
a = 8'd144; b = 8'd190;  #10 
a = 8'd144; b = 8'd191;  #10 
a = 8'd144; b = 8'd192;  #10 
a = 8'd144; b = 8'd193;  #10 
a = 8'd144; b = 8'd194;  #10 
a = 8'd144; b = 8'd195;  #10 
a = 8'd144; b = 8'd196;  #10 
a = 8'd144; b = 8'd197;  #10 
a = 8'd144; b = 8'd198;  #10 
a = 8'd144; b = 8'd199;  #10 
a = 8'd144; b = 8'd200;  #10 
a = 8'd144; b = 8'd201;  #10 
a = 8'd144; b = 8'd202;  #10 
a = 8'd144; b = 8'd203;  #10 
a = 8'd144; b = 8'd204;  #10 
a = 8'd144; b = 8'd205;  #10 
a = 8'd144; b = 8'd206;  #10 
a = 8'd144; b = 8'd207;  #10 
a = 8'd144; b = 8'd208;  #10 
a = 8'd144; b = 8'd209;  #10 
a = 8'd144; b = 8'd210;  #10 
a = 8'd144; b = 8'd211;  #10 
a = 8'd144; b = 8'd212;  #10 
a = 8'd144; b = 8'd213;  #10 
a = 8'd144; b = 8'd214;  #10 
a = 8'd144; b = 8'd215;  #10 
a = 8'd144; b = 8'd216;  #10 
a = 8'd144; b = 8'd217;  #10 
a = 8'd144; b = 8'd218;  #10 
a = 8'd144; b = 8'd219;  #10 
a = 8'd144; b = 8'd220;  #10 
a = 8'd144; b = 8'd221;  #10 
a = 8'd144; b = 8'd222;  #10 
a = 8'd144; b = 8'd223;  #10 
a = 8'd144; b = 8'd224;  #10 
a = 8'd144; b = 8'd225;  #10 
a = 8'd144; b = 8'd226;  #10 
a = 8'd144; b = 8'd227;  #10 
a = 8'd144; b = 8'd228;  #10 
a = 8'd144; b = 8'd229;  #10 
a = 8'd144; b = 8'd230;  #10 
a = 8'd144; b = 8'd231;  #10 
a = 8'd144; b = 8'd232;  #10 
a = 8'd144; b = 8'd233;  #10 
a = 8'd144; b = 8'd234;  #10 
a = 8'd144; b = 8'd235;  #10 
a = 8'd144; b = 8'd236;  #10 
a = 8'd144; b = 8'd237;  #10 
a = 8'd144; b = 8'd238;  #10 
a = 8'd144; b = 8'd239;  #10 
a = 8'd144; b = 8'd240;  #10 
a = 8'd144; b = 8'd241;  #10 
a = 8'd144; b = 8'd242;  #10 
a = 8'd144; b = 8'd243;  #10 
a = 8'd144; b = 8'd244;  #10 
a = 8'd144; b = 8'd245;  #10 
a = 8'd144; b = 8'd246;  #10 
a = 8'd144; b = 8'd247;  #10 
a = 8'd144; b = 8'd248;  #10 
a = 8'd144; b = 8'd249;  #10 
a = 8'd144; b = 8'd250;  #10 
a = 8'd144; b = 8'd251;  #10 
a = 8'd144; b = 8'd252;  #10 
a = 8'd144; b = 8'd253;  #10 
a = 8'd144; b = 8'd254;  #10 
a = 8'd144; b = 8'd255;  #10 
a = 8'd145; b = 8'd0;  #10 
a = 8'd145; b = 8'd1;  #10 
a = 8'd145; b = 8'd2;  #10 
a = 8'd145; b = 8'd3;  #10 
a = 8'd145; b = 8'd4;  #10 
a = 8'd145; b = 8'd5;  #10 
a = 8'd145; b = 8'd6;  #10 
a = 8'd145; b = 8'd7;  #10 
a = 8'd145; b = 8'd8;  #10 
a = 8'd145; b = 8'd9;  #10 
a = 8'd145; b = 8'd10;  #10 
a = 8'd145; b = 8'd11;  #10 
a = 8'd145; b = 8'd12;  #10 
a = 8'd145; b = 8'd13;  #10 
a = 8'd145; b = 8'd14;  #10 
a = 8'd145; b = 8'd15;  #10 
a = 8'd145; b = 8'd16;  #10 
a = 8'd145; b = 8'd17;  #10 
a = 8'd145; b = 8'd18;  #10 
a = 8'd145; b = 8'd19;  #10 
a = 8'd145; b = 8'd20;  #10 
a = 8'd145; b = 8'd21;  #10 
a = 8'd145; b = 8'd22;  #10 
a = 8'd145; b = 8'd23;  #10 
a = 8'd145; b = 8'd24;  #10 
a = 8'd145; b = 8'd25;  #10 
a = 8'd145; b = 8'd26;  #10 
a = 8'd145; b = 8'd27;  #10 
a = 8'd145; b = 8'd28;  #10 
a = 8'd145; b = 8'd29;  #10 
a = 8'd145; b = 8'd30;  #10 
a = 8'd145; b = 8'd31;  #10 
a = 8'd145; b = 8'd32;  #10 
a = 8'd145; b = 8'd33;  #10 
a = 8'd145; b = 8'd34;  #10 
a = 8'd145; b = 8'd35;  #10 
a = 8'd145; b = 8'd36;  #10 
a = 8'd145; b = 8'd37;  #10 
a = 8'd145; b = 8'd38;  #10 
a = 8'd145; b = 8'd39;  #10 
a = 8'd145; b = 8'd40;  #10 
a = 8'd145; b = 8'd41;  #10 
a = 8'd145; b = 8'd42;  #10 
a = 8'd145; b = 8'd43;  #10 
a = 8'd145; b = 8'd44;  #10 
a = 8'd145; b = 8'd45;  #10 
a = 8'd145; b = 8'd46;  #10 
a = 8'd145; b = 8'd47;  #10 
a = 8'd145; b = 8'd48;  #10 
a = 8'd145; b = 8'd49;  #10 
a = 8'd145; b = 8'd50;  #10 
a = 8'd145; b = 8'd51;  #10 
a = 8'd145; b = 8'd52;  #10 
a = 8'd145; b = 8'd53;  #10 
a = 8'd145; b = 8'd54;  #10 
a = 8'd145; b = 8'd55;  #10 
a = 8'd145; b = 8'd56;  #10 
a = 8'd145; b = 8'd57;  #10 
a = 8'd145; b = 8'd58;  #10 
a = 8'd145; b = 8'd59;  #10 
a = 8'd145; b = 8'd60;  #10 
a = 8'd145; b = 8'd61;  #10 
a = 8'd145; b = 8'd62;  #10 
a = 8'd145; b = 8'd63;  #10 
a = 8'd145; b = 8'd64;  #10 
a = 8'd145; b = 8'd65;  #10 
a = 8'd145; b = 8'd66;  #10 
a = 8'd145; b = 8'd67;  #10 
a = 8'd145; b = 8'd68;  #10 
a = 8'd145; b = 8'd69;  #10 
a = 8'd145; b = 8'd70;  #10 
a = 8'd145; b = 8'd71;  #10 
a = 8'd145; b = 8'd72;  #10 
a = 8'd145; b = 8'd73;  #10 
a = 8'd145; b = 8'd74;  #10 
a = 8'd145; b = 8'd75;  #10 
a = 8'd145; b = 8'd76;  #10 
a = 8'd145; b = 8'd77;  #10 
a = 8'd145; b = 8'd78;  #10 
a = 8'd145; b = 8'd79;  #10 
a = 8'd145; b = 8'd80;  #10 
a = 8'd145; b = 8'd81;  #10 
a = 8'd145; b = 8'd82;  #10 
a = 8'd145; b = 8'd83;  #10 
a = 8'd145; b = 8'd84;  #10 
a = 8'd145; b = 8'd85;  #10 
a = 8'd145; b = 8'd86;  #10 
a = 8'd145; b = 8'd87;  #10 
a = 8'd145; b = 8'd88;  #10 
a = 8'd145; b = 8'd89;  #10 
a = 8'd145; b = 8'd90;  #10 
a = 8'd145; b = 8'd91;  #10 
a = 8'd145; b = 8'd92;  #10 
a = 8'd145; b = 8'd93;  #10 
a = 8'd145; b = 8'd94;  #10 
a = 8'd145; b = 8'd95;  #10 
a = 8'd145; b = 8'd96;  #10 
a = 8'd145; b = 8'd97;  #10 
a = 8'd145; b = 8'd98;  #10 
a = 8'd145; b = 8'd99;  #10 
a = 8'd145; b = 8'd100;  #10 
a = 8'd145; b = 8'd101;  #10 
a = 8'd145; b = 8'd102;  #10 
a = 8'd145; b = 8'd103;  #10 
a = 8'd145; b = 8'd104;  #10 
a = 8'd145; b = 8'd105;  #10 
a = 8'd145; b = 8'd106;  #10 
a = 8'd145; b = 8'd107;  #10 
a = 8'd145; b = 8'd108;  #10 
a = 8'd145; b = 8'd109;  #10 
a = 8'd145; b = 8'd110;  #10 
a = 8'd145; b = 8'd111;  #10 
a = 8'd145; b = 8'd112;  #10 
a = 8'd145; b = 8'd113;  #10 
a = 8'd145; b = 8'd114;  #10 
a = 8'd145; b = 8'd115;  #10 
a = 8'd145; b = 8'd116;  #10 
a = 8'd145; b = 8'd117;  #10 
a = 8'd145; b = 8'd118;  #10 
a = 8'd145; b = 8'd119;  #10 
a = 8'd145; b = 8'd120;  #10 
a = 8'd145; b = 8'd121;  #10 
a = 8'd145; b = 8'd122;  #10 
a = 8'd145; b = 8'd123;  #10 
a = 8'd145; b = 8'd124;  #10 
a = 8'd145; b = 8'd125;  #10 
a = 8'd145; b = 8'd126;  #10 
a = 8'd145; b = 8'd127;  #10 
a = 8'd145; b = 8'd128;  #10 
a = 8'd145; b = 8'd129;  #10 
a = 8'd145; b = 8'd130;  #10 
a = 8'd145; b = 8'd131;  #10 
a = 8'd145; b = 8'd132;  #10 
a = 8'd145; b = 8'd133;  #10 
a = 8'd145; b = 8'd134;  #10 
a = 8'd145; b = 8'd135;  #10 
a = 8'd145; b = 8'd136;  #10 
a = 8'd145; b = 8'd137;  #10 
a = 8'd145; b = 8'd138;  #10 
a = 8'd145; b = 8'd139;  #10 
a = 8'd145; b = 8'd140;  #10 
a = 8'd145; b = 8'd141;  #10 
a = 8'd145; b = 8'd142;  #10 
a = 8'd145; b = 8'd143;  #10 
a = 8'd145; b = 8'd144;  #10 
a = 8'd145; b = 8'd145;  #10 
a = 8'd145; b = 8'd146;  #10 
a = 8'd145; b = 8'd147;  #10 
a = 8'd145; b = 8'd148;  #10 
a = 8'd145; b = 8'd149;  #10 
a = 8'd145; b = 8'd150;  #10 
a = 8'd145; b = 8'd151;  #10 
a = 8'd145; b = 8'd152;  #10 
a = 8'd145; b = 8'd153;  #10 
a = 8'd145; b = 8'd154;  #10 
a = 8'd145; b = 8'd155;  #10 
a = 8'd145; b = 8'd156;  #10 
a = 8'd145; b = 8'd157;  #10 
a = 8'd145; b = 8'd158;  #10 
a = 8'd145; b = 8'd159;  #10 
a = 8'd145; b = 8'd160;  #10 
a = 8'd145; b = 8'd161;  #10 
a = 8'd145; b = 8'd162;  #10 
a = 8'd145; b = 8'd163;  #10 
a = 8'd145; b = 8'd164;  #10 
a = 8'd145; b = 8'd165;  #10 
a = 8'd145; b = 8'd166;  #10 
a = 8'd145; b = 8'd167;  #10 
a = 8'd145; b = 8'd168;  #10 
a = 8'd145; b = 8'd169;  #10 
a = 8'd145; b = 8'd170;  #10 
a = 8'd145; b = 8'd171;  #10 
a = 8'd145; b = 8'd172;  #10 
a = 8'd145; b = 8'd173;  #10 
a = 8'd145; b = 8'd174;  #10 
a = 8'd145; b = 8'd175;  #10 
a = 8'd145; b = 8'd176;  #10 
a = 8'd145; b = 8'd177;  #10 
a = 8'd145; b = 8'd178;  #10 
a = 8'd145; b = 8'd179;  #10 
a = 8'd145; b = 8'd180;  #10 
a = 8'd145; b = 8'd181;  #10 
a = 8'd145; b = 8'd182;  #10 
a = 8'd145; b = 8'd183;  #10 
a = 8'd145; b = 8'd184;  #10 
a = 8'd145; b = 8'd185;  #10 
a = 8'd145; b = 8'd186;  #10 
a = 8'd145; b = 8'd187;  #10 
a = 8'd145; b = 8'd188;  #10 
a = 8'd145; b = 8'd189;  #10 
a = 8'd145; b = 8'd190;  #10 
a = 8'd145; b = 8'd191;  #10 
a = 8'd145; b = 8'd192;  #10 
a = 8'd145; b = 8'd193;  #10 
a = 8'd145; b = 8'd194;  #10 
a = 8'd145; b = 8'd195;  #10 
a = 8'd145; b = 8'd196;  #10 
a = 8'd145; b = 8'd197;  #10 
a = 8'd145; b = 8'd198;  #10 
a = 8'd145; b = 8'd199;  #10 
a = 8'd145; b = 8'd200;  #10 
a = 8'd145; b = 8'd201;  #10 
a = 8'd145; b = 8'd202;  #10 
a = 8'd145; b = 8'd203;  #10 
a = 8'd145; b = 8'd204;  #10 
a = 8'd145; b = 8'd205;  #10 
a = 8'd145; b = 8'd206;  #10 
a = 8'd145; b = 8'd207;  #10 
a = 8'd145; b = 8'd208;  #10 
a = 8'd145; b = 8'd209;  #10 
a = 8'd145; b = 8'd210;  #10 
a = 8'd145; b = 8'd211;  #10 
a = 8'd145; b = 8'd212;  #10 
a = 8'd145; b = 8'd213;  #10 
a = 8'd145; b = 8'd214;  #10 
a = 8'd145; b = 8'd215;  #10 
a = 8'd145; b = 8'd216;  #10 
a = 8'd145; b = 8'd217;  #10 
a = 8'd145; b = 8'd218;  #10 
a = 8'd145; b = 8'd219;  #10 
a = 8'd145; b = 8'd220;  #10 
a = 8'd145; b = 8'd221;  #10 
a = 8'd145; b = 8'd222;  #10 
a = 8'd145; b = 8'd223;  #10 
a = 8'd145; b = 8'd224;  #10 
a = 8'd145; b = 8'd225;  #10 
a = 8'd145; b = 8'd226;  #10 
a = 8'd145; b = 8'd227;  #10 
a = 8'd145; b = 8'd228;  #10 
a = 8'd145; b = 8'd229;  #10 
a = 8'd145; b = 8'd230;  #10 
a = 8'd145; b = 8'd231;  #10 
a = 8'd145; b = 8'd232;  #10 
a = 8'd145; b = 8'd233;  #10 
a = 8'd145; b = 8'd234;  #10 
a = 8'd145; b = 8'd235;  #10 
a = 8'd145; b = 8'd236;  #10 
a = 8'd145; b = 8'd237;  #10 
a = 8'd145; b = 8'd238;  #10 
a = 8'd145; b = 8'd239;  #10 
a = 8'd145; b = 8'd240;  #10 
a = 8'd145; b = 8'd241;  #10 
a = 8'd145; b = 8'd242;  #10 
a = 8'd145; b = 8'd243;  #10 
a = 8'd145; b = 8'd244;  #10 
a = 8'd145; b = 8'd245;  #10 
a = 8'd145; b = 8'd246;  #10 
a = 8'd145; b = 8'd247;  #10 
a = 8'd145; b = 8'd248;  #10 
a = 8'd145; b = 8'd249;  #10 
a = 8'd145; b = 8'd250;  #10 
a = 8'd145; b = 8'd251;  #10 
a = 8'd145; b = 8'd252;  #10 
a = 8'd145; b = 8'd253;  #10 
a = 8'd145; b = 8'd254;  #10 
a = 8'd145; b = 8'd255;  #10 
a = 8'd146; b = 8'd0;  #10 
a = 8'd146; b = 8'd1;  #10 
a = 8'd146; b = 8'd2;  #10 
a = 8'd146; b = 8'd3;  #10 
a = 8'd146; b = 8'd4;  #10 
a = 8'd146; b = 8'd5;  #10 
a = 8'd146; b = 8'd6;  #10 
a = 8'd146; b = 8'd7;  #10 
a = 8'd146; b = 8'd8;  #10 
a = 8'd146; b = 8'd9;  #10 
a = 8'd146; b = 8'd10;  #10 
a = 8'd146; b = 8'd11;  #10 
a = 8'd146; b = 8'd12;  #10 
a = 8'd146; b = 8'd13;  #10 
a = 8'd146; b = 8'd14;  #10 
a = 8'd146; b = 8'd15;  #10 
a = 8'd146; b = 8'd16;  #10 
a = 8'd146; b = 8'd17;  #10 
a = 8'd146; b = 8'd18;  #10 
a = 8'd146; b = 8'd19;  #10 
a = 8'd146; b = 8'd20;  #10 
a = 8'd146; b = 8'd21;  #10 
a = 8'd146; b = 8'd22;  #10 
a = 8'd146; b = 8'd23;  #10 
a = 8'd146; b = 8'd24;  #10 
a = 8'd146; b = 8'd25;  #10 
a = 8'd146; b = 8'd26;  #10 
a = 8'd146; b = 8'd27;  #10 
a = 8'd146; b = 8'd28;  #10 
a = 8'd146; b = 8'd29;  #10 
a = 8'd146; b = 8'd30;  #10 
a = 8'd146; b = 8'd31;  #10 
a = 8'd146; b = 8'd32;  #10 
a = 8'd146; b = 8'd33;  #10 
a = 8'd146; b = 8'd34;  #10 
a = 8'd146; b = 8'd35;  #10 
a = 8'd146; b = 8'd36;  #10 
a = 8'd146; b = 8'd37;  #10 
a = 8'd146; b = 8'd38;  #10 
a = 8'd146; b = 8'd39;  #10 
a = 8'd146; b = 8'd40;  #10 
a = 8'd146; b = 8'd41;  #10 
a = 8'd146; b = 8'd42;  #10 
a = 8'd146; b = 8'd43;  #10 
a = 8'd146; b = 8'd44;  #10 
a = 8'd146; b = 8'd45;  #10 
a = 8'd146; b = 8'd46;  #10 
a = 8'd146; b = 8'd47;  #10 
a = 8'd146; b = 8'd48;  #10 
a = 8'd146; b = 8'd49;  #10 
a = 8'd146; b = 8'd50;  #10 
a = 8'd146; b = 8'd51;  #10 
a = 8'd146; b = 8'd52;  #10 
a = 8'd146; b = 8'd53;  #10 
a = 8'd146; b = 8'd54;  #10 
a = 8'd146; b = 8'd55;  #10 
a = 8'd146; b = 8'd56;  #10 
a = 8'd146; b = 8'd57;  #10 
a = 8'd146; b = 8'd58;  #10 
a = 8'd146; b = 8'd59;  #10 
a = 8'd146; b = 8'd60;  #10 
a = 8'd146; b = 8'd61;  #10 
a = 8'd146; b = 8'd62;  #10 
a = 8'd146; b = 8'd63;  #10 
a = 8'd146; b = 8'd64;  #10 
a = 8'd146; b = 8'd65;  #10 
a = 8'd146; b = 8'd66;  #10 
a = 8'd146; b = 8'd67;  #10 
a = 8'd146; b = 8'd68;  #10 
a = 8'd146; b = 8'd69;  #10 
a = 8'd146; b = 8'd70;  #10 
a = 8'd146; b = 8'd71;  #10 
a = 8'd146; b = 8'd72;  #10 
a = 8'd146; b = 8'd73;  #10 
a = 8'd146; b = 8'd74;  #10 
a = 8'd146; b = 8'd75;  #10 
a = 8'd146; b = 8'd76;  #10 
a = 8'd146; b = 8'd77;  #10 
a = 8'd146; b = 8'd78;  #10 
a = 8'd146; b = 8'd79;  #10 
a = 8'd146; b = 8'd80;  #10 
a = 8'd146; b = 8'd81;  #10 
a = 8'd146; b = 8'd82;  #10 
a = 8'd146; b = 8'd83;  #10 
a = 8'd146; b = 8'd84;  #10 
a = 8'd146; b = 8'd85;  #10 
a = 8'd146; b = 8'd86;  #10 
a = 8'd146; b = 8'd87;  #10 
a = 8'd146; b = 8'd88;  #10 
a = 8'd146; b = 8'd89;  #10 
a = 8'd146; b = 8'd90;  #10 
a = 8'd146; b = 8'd91;  #10 
a = 8'd146; b = 8'd92;  #10 
a = 8'd146; b = 8'd93;  #10 
a = 8'd146; b = 8'd94;  #10 
a = 8'd146; b = 8'd95;  #10 
a = 8'd146; b = 8'd96;  #10 
a = 8'd146; b = 8'd97;  #10 
a = 8'd146; b = 8'd98;  #10 
a = 8'd146; b = 8'd99;  #10 
a = 8'd146; b = 8'd100;  #10 
a = 8'd146; b = 8'd101;  #10 
a = 8'd146; b = 8'd102;  #10 
a = 8'd146; b = 8'd103;  #10 
a = 8'd146; b = 8'd104;  #10 
a = 8'd146; b = 8'd105;  #10 
a = 8'd146; b = 8'd106;  #10 
a = 8'd146; b = 8'd107;  #10 
a = 8'd146; b = 8'd108;  #10 
a = 8'd146; b = 8'd109;  #10 
a = 8'd146; b = 8'd110;  #10 
a = 8'd146; b = 8'd111;  #10 
a = 8'd146; b = 8'd112;  #10 
a = 8'd146; b = 8'd113;  #10 
a = 8'd146; b = 8'd114;  #10 
a = 8'd146; b = 8'd115;  #10 
a = 8'd146; b = 8'd116;  #10 
a = 8'd146; b = 8'd117;  #10 
a = 8'd146; b = 8'd118;  #10 
a = 8'd146; b = 8'd119;  #10 
a = 8'd146; b = 8'd120;  #10 
a = 8'd146; b = 8'd121;  #10 
a = 8'd146; b = 8'd122;  #10 
a = 8'd146; b = 8'd123;  #10 
a = 8'd146; b = 8'd124;  #10 
a = 8'd146; b = 8'd125;  #10 
a = 8'd146; b = 8'd126;  #10 
a = 8'd146; b = 8'd127;  #10 
a = 8'd146; b = 8'd128;  #10 
a = 8'd146; b = 8'd129;  #10 
a = 8'd146; b = 8'd130;  #10 
a = 8'd146; b = 8'd131;  #10 
a = 8'd146; b = 8'd132;  #10 
a = 8'd146; b = 8'd133;  #10 
a = 8'd146; b = 8'd134;  #10 
a = 8'd146; b = 8'd135;  #10 
a = 8'd146; b = 8'd136;  #10 
a = 8'd146; b = 8'd137;  #10 
a = 8'd146; b = 8'd138;  #10 
a = 8'd146; b = 8'd139;  #10 
a = 8'd146; b = 8'd140;  #10 
a = 8'd146; b = 8'd141;  #10 
a = 8'd146; b = 8'd142;  #10 
a = 8'd146; b = 8'd143;  #10 
a = 8'd146; b = 8'd144;  #10 
a = 8'd146; b = 8'd145;  #10 
a = 8'd146; b = 8'd146;  #10 
a = 8'd146; b = 8'd147;  #10 
a = 8'd146; b = 8'd148;  #10 
a = 8'd146; b = 8'd149;  #10 
a = 8'd146; b = 8'd150;  #10 
a = 8'd146; b = 8'd151;  #10 
a = 8'd146; b = 8'd152;  #10 
a = 8'd146; b = 8'd153;  #10 
a = 8'd146; b = 8'd154;  #10 
a = 8'd146; b = 8'd155;  #10 
a = 8'd146; b = 8'd156;  #10 
a = 8'd146; b = 8'd157;  #10 
a = 8'd146; b = 8'd158;  #10 
a = 8'd146; b = 8'd159;  #10 
a = 8'd146; b = 8'd160;  #10 
a = 8'd146; b = 8'd161;  #10 
a = 8'd146; b = 8'd162;  #10 
a = 8'd146; b = 8'd163;  #10 
a = 8'd146; b = 8'd164;  #10 
a = 8'd146; b = 8'd165;  #10 
a = 8'd146; b = 8'd166;  #10 
a = 8'd146; b = 8'd167;  #10 
a = 8'd146; b = 8'd168;  #10 
a = 8'd146; b = 8'd169;  #10 
a = 8'd146; b = 8'd170;  #10 
a = 8'd146; b = 8'd171;  #10 
a = 8'd146; b = 8'd172;  #10 
a = 8'd146; b = 8'd173;  #10 
a = 8'd146; b = 8'd174;  #10 
a = 8'd146; b = 8'd175;  #10 
a = 8'd146; b = 8'd176;  #10 
a = 8'd146; b = 8'd177;  #10 
a = 8'd146; b = 8'd178;  #10 
a = 8'd146; b = 8'd179;  #10 
a = 8'd146; b = 8'd180;  #10 
a = 8'd146; b = 8'd181;  #10 
a = 8'd146; b = 8'd182;  #10 
a = 8'd146; b = 8'd183;  #10 
a = 8'd146; b = 8'd184;  #10 
a = 8'd146; b = 8'd185;  #10 
a = 8'd146; b = 8'd186;  #10 
a = 8'd146; b = 8'd187;  #10 
a = 8'd146; b = 8'd188;  #10 
a = 8'd146; b = 8'd189;  #10 
a = 8'd146; b = 8'd190;  #10 
a = 8'd146; b = 8'd191;  #10 
a = 8'd146; b = 8'd192;  #10 
a = 8'd146; b = 8'd193;  #10 
a = 8'd146; b = 8'd194;  #10 
a = 8'd146; b = 8'd195;  #10 
a = 8'd146; b = 8'd196;  #10 
a = 8'd146; b = 8'd197;  #10 
a = 8'd146; b = 8'd198;  #10 
a = 8'd146; b = 8'd199;  #10 
a = 8'd146; b = 8'd200;  #10 
a = 8'd146; b = 8'd201;  #10 
a = 8'd146; b = 8'd202;  #10 
a = 8'd146; b = 8'd203;  #10 
a = 8'd146; b = 8'd204;  #10 
a = 8'd146; b = 8'd205;  #10 
a = 8'd146; b = 8'd206;  #10 
a = 8'd146; b = 8'd207;  #10 
a = 8'd146; b = 8'd208;  #10 
a = 8'd146; b = 8'd209;  #10 
a = 8'd146; b = 8'd210;  #10 
a = 8'd146; b = 8'd211;  #10 
a = 8'd146; b = 8'd212;  #10 
a = 8'd146; b = 8'd213;  #10 
a = 8'd146; b = 8'd214;  #10 
a = 8'd146; b = 8'd215;  #10 
a = 8'd146; b = 8'd216;  #10 
a = 8'd146; b = 8'd217;  #10 
a = 8'd146; b = 8'd218;  #10 
a = 8'd146; b = 8'd219;  #10 
a = 8'd146; b = 8'd220;  #10 
a = 8'd146; b = 8'd221;  #10 
a = 8'd146; b = 8'd222;  #10 
a = 8'd146; b = 8'd223;  #10 
a = 8'd146; b = 8'd224;  #10 
a = 8'd146; b = 8'd225;  #10 
a = 8'd146; b = 8'd226;  #10 
a = 8'd146; b = 8'd227;  #10 
a = 8'd146; b = 8'd228;  #10 
a = 8'd146; b = 8'd229;  #10 
a = 8'd146; b = 8'd230;  #10 
a = 8'd146; b = 8'd231;  #10 
a = 8'd146; b = 8'd232;  #10 
a = 8'd146; b = 8'd233;  #10 
a = 8'd146; b = 8'd234;  #10 
a = 8'd146; b = 8'd235;  #10 
a = 8'd146; b = 8'd236;  #10 
a = 8'd146; b = 8'd237;  #10 
a = 8'd146; b = 8'd238;  #10 
a = 8'd146; b = 8'd239;  #10 
a = 8'd146; b = 8'd240;  #10 
a = 8'd146; b = 8'd241;  #10 
a = 8'd146; b = 8'd242;  #10 
a = 8'd146; b = 8'd243;  #10 
a = 8'd146; b = 8'd244;  #10 
a = 8'd146; b = 8'd245;  #10 
a = 8'd146; b = 8'd246;  #10 
a = 8'd146; b = 8'd247;  #10 
a = 8'd146; b = 8'd248;  #10 
a = 8'd146; b = 8'd249;  #10 
a = 8'd146; b = 8'd250;  #10 
a = 8'd146; b = 8'd251;  #10 
a = 8'd146; b = 8'd252;  #10 
a = 8'd146; b = 8'd253;  #10 
a = 8'd146; b = 8'd254;  #10 
a = 8'd146; b = 8'd255;  #10 
a = 8'd147; b = 8'd0;  #10 
a = 8'd147; b = 8'd1;  #10 
a = 8'd147; b = 8'd2;  #10 
a = 8'd147; b = 8'd3;  #10 
a = 8'd147; b = 8'd4;  #10 
a = 8'd147; b = 8'd5;  #10 
a = 8'd147; b = 8'd6;  #10 
a = 8'd147; b = 8'd7;  #10 
a = 8'd147; b = 8'd8;  #10 
a = 8'd147; b = 8'd9;  #10 
a = 8'd147; b = 8'd10;  #10 
a = 8'd147; b = 8'd11;  #10 
a = 8'd147; b = 8'd12;  #10 
a = 8'd147; b = 8'd13;  #10 
a = 8'd147; b = 8'd14;  #10 
a = 8'd147; b = 8'd15;  #10 
a = 8'd147; b = 8'd16;  #10 
a = 8'd147; b = 8'd17;  #10 
a = 8'd147; b = 8'd18;  #10 
a = 8'd147; b = 8'd19;  #10 
a = 8'd147; b = 8'd20;  #10 
a = 8'd147; b = 8'd21;  #10 
a = 8'd147; b = 8'd22;  #10 
a = 8'd147; b = 8'd23;  #10 
a = 8'd147; b = 8'd24;  #10 
a = 8'd147; b = 8'd25;  #10 
a = 8'd147; b = 8'd26;  #10 
a = 8'd147; b = 8'd27;  #10 
a = 8'd147; b = 8'd28;  #10 
a = 8'd147; b = 8'd29;  #10 
a = 8'd147; b = 8'd30;  #10 
a = 8'd147; b = 8'd31;  #10 
a = 8'd147; b = 8'd32;  #10 
a = 8'd147; b = 8'd33;  #10 
a = 8'd147; b = 8'd34;  #10 
a = 8'd147; b = 8'd35;  #10 
a = 8'd147; b = 8'd36;  #10 
a = 8'd147; b = 8'd37;  #10 
a = 8'd147; b = 8'd38;  #10 
a = 8'd147; b = 8'd39;  #10 
a = 8'd147; b = 8'd40;  #10 
a = 8'd147; b = 8'd41;  #10 
a = 8'd147; b = 8'd42;  #10 
a = 8'd147; b = 8'd43;  #10 
a = 8'd147; b = 8'd44;  #10 
a = 8'd147; b = 8'd45;  #10 
a = 8'd147; b = 8'd46;  #10 
a = 8'd147; b = 8'd47;  #10 
a = 8'd147; b = 8'd48;  #10 
a = 8'd147; b = 8'd49;  #10 
a = 8'd147; b = 8'd50;  #10 
a = 8'd147; b = 8'd51;  #10 
a = 8'd147; b = 8'd52;  #10 
a = 8'd147; b = 8'd53;  #10 
a = 8'd147; b = 8'd54;  #10 
a = 8'd147; b = 8'd55;  #10 
a = 8'd147; b = 8'd56;  #10 
a = 8'd147; b = 8'd57;  #10 
a = 8'd147; b = 8'd58;  #10 
a = 8'd147; b = 8'd59;  #10 
a = 8'd147; b = 8'd60;  #10 
a = 8'd147; b = 8'd61;  #10 
a = 8'd147; b = 8'd62;  #10 
a = 8'd147; b = 8'd63;  #10 
a = 8'd147; b = 8'd64;  #10 
a = 8'd147; b = 8'd65;  #10 
a = 8'd147; b = 8'd66;  #10 
a = 8'd147; b = 8'd67;  #10 
a = 8'd147; b = 8'd68;  #10 
a = 8'd147; b = 8'd69;  #10 
a = 8'd147; b = 8'd70;  #10 
a = 8'd147; b = 8'd71;  #10 
a = 8'd147; b = 8'd72;  #10 
a = 8'd147; b = 8'd73;  #10 
a = 8'd147; b = 8'd74;  #10 
a = 8'd147; b = 8'd75;  #10 
a = 8'd147; b = 8'd76;  #10 
a = 8'd147; b = 8'd77;  #10 
a = 8'd147; b = 8'd78;  #10 
a = 8'd147; b = 8'd79;  #10 
a = 8'd147; b = 8'd80;  #10 
a = 8'd147; b = 8'd81;  #10 
a = 8'd147; b = 8'd82;  #10 
a = 8'd147; b = 8'd83;  #10 
a = 8'd147; b = 8'd84;  #10 
a = 8'd147; b = 8'd85;  #10 
a = 8'd147; b = 8'd86;  #10 
a = 8'd147; b = 8'd87;  #10 
a = 8'd147; b = 8'd88;  #10 
a = 8'd147; b = 8'd89;  #10 
a = 8'd147; b = 8'd90;  #10 
a = 8'd147; b = 8'd91;  #10 
a = 8'd147; b = 8'd92;  #10 
a = 8'd147; b = 8'd93;  #10 
a = 8'd147; b = 8'd94;  #10 
a = 8'd147; b = 8'd95;  #10 
a = 8'd147; b = 8'd96;  #10 
a = 8'd147; b = 8'd97;  #10 
a = 8'd147; b = 8'd98;  #10 
a = 8'd147; b = 8'd99;  #10 
a = 8'd147; b = 8'd100;  #10 
a = 8'd147; b = 8'd101;  #10 
a = 8'd147; b = 8'd102;  #10 
a = 8'd147; b = 8'd103;  #10 
a = 8'd147; b = 8'd104;  #10 
a = 8'd147; b = 8'd105;  #10 
a = 8'd147; b = 8'd106;  #10 
a = 8'd147; b = 8'd107;  #10 
a = 8'd147; b = 8'd108;  #10 
a = 8'd147; b = 8'd109;  #10 
a = 8'd147; b = 8'd110;  #10 
a = 8'd147; b = 8'd111;  #10 
a = 8'd147; b = 8'd112;  #10 
a = 8'd147; b = 8'd113;  #10 
a = 8'd147; b = 8'd114;  #10 
a = 8'd147; b = 8'd115;  #10 
a = 8'd147; b = 8'd116;  #10 
a = 8'd147; b = 8'd117;  #10 
a = 8'd147; b = 8'd118;  #10 
a = 8'd147; b = 8'd119;  #10 
a = 8'd147; b = 8'd120;  #10 
a = 8'd147; b = 8'd121;  #10 
a = 8'd147; b = 8'd122;  #10 
a = 8'd147; b = 8'd123;  #10 
a = 8'd147; b = 8'd124;  #10 
a = 8'd147; b = 8'd125;  #10 
a = 8'd147; b = 8'd126;  #10 
a = 8'd147; b = 8'd127;  #10 
a = 8'd147; b = 8'd128;  #10 
a = 8'd147; b = 8'd129;  #10 
a = 8'd147; b = 8'd130;  #10 
a = 8'd147; b = 8'd131;  #10 
a = 8'd147; b = 8'd132;  #10 
a = 8'd147; b = 8'd133;  #10 
a = 8'd147; b = 8'd134;  #10 
a = 8'd147; b = 8'd135;  #10 
a = 8'd147; b = 8'd136;  #10 
a = 8'd147; b = 8'd137;  #10 
a = 8'd147; b = 8'd138;  #10 
a = 8'd147; b = 8'd139;  #10 
a = 8'd147; b = 8'd140;  #10 
a = 8'd147; b = 8'd141;  #10 
a = 8'd147; b = 8'd142;  #10 
a = 8'd147; b = 8'd143;  #10 
a = 8'd147; b = 8'd144;  #10 
a = 8'd147; b = 8'd145;  #10 
a = 8'd147; b = 8'd146;  #10 
a = 8'd147; b = 8'd147;  #10 
a = 8'd147; b = 8'd148;  #10 
a = 8'd147; b = 8'd149;  #10 
a = 8'd147; b = 8'd150;  #10 
a = 8'd147; b = 8'd151;  #10 
a = 8'd147; b = 8'd152;  #10 
a = 8'd147; b = 8'd153;  #10 
a = 8'd147; b = 8'd154;  #10 
a = 8'd147; b = 8'd155;  #10 
a = 8'd147; b = 8'd156;  #10 
a = 8'd147; b = 8'd157;  #10 
a = 8'd147; b = 8'd158;  #10 
a = 8'd147; b = 8'd159;  #10 
a = 8'd147; b = 8'd160;  #10 
a = 8'd147; b = 8'd161;  #10 
a = 8'd147; b = 8'd162;  #10 
a = 8'd147; b = 8'd163;  #10 
a = 8'd147; b = 8'd164;  #10 
a = 8'd147; b = 8'd165;  #10 
a = 8'd147; b = 8'd166;  #10 
a = 8'd147; b = 8'd167;  #10 
a = 8'd147; b = 8'd168;  #10 
a = 8'd147; b = 8'd169;  #10 
a = 8'd147; b = 8'd170;  #10 
a = 8'd147; b = 8'd171;  #10 
a = 8'd147; b = 8'd172;  #10 
a = 8'd147; b = 8'd173;  #10 
a = 8'd147; b = 8'd174;  #10 
a = 8'd147; b = 8'd175;  #10 
a = 8'd147; b = 8'd176;  #10 
a = 8'd147; b = 8'd177;  #10 
a = 8'd147; b = 8'd178;  #10 
a = 8'd147; b = 8'd179;  #10 
a = 8'd147; b = 8'd180;  #10 
a = 8'd147; b = 8'd181;  #10 
a = 8'd147; b = 8'd182;  #10 
a = 8'd147; b = 8'd183;  #10 
a = 8'd147; b = 8'd184;  #10 
a = 8'd147; b = 8'd185;  #10 
a = 8'd147; b = 8'd186;  #10 
a = 8'd147; b = 8'd187;  #10 
a = 8'd147; b = 8'd188;  #10 
a = 8'd147; b = 8'd189;  #10 
a = 8'd147; b = 8'd190;  #10 
a = 8'd147; b = 8'd191;  #10 
a = 8'd147; b = 8'd192;  #10 
a = 8'd147; b = 8'd193;  #10 
a = 8'd147; b = 8'd194;  #10 
a = 8'd147; b = 8'd195;  #10 
a = 8'd147; b = 8'd196;  #10 
a = 8'd147; b = 8'd197;  #10 
a = 8'd147; b = 8'd198;  #10 
a = 8'd147; b = 8'd199;  #10 
a = 8'd147; b = 8'd200;  #10 
a = 8'd147; b = 8'd201;  #10 
a = 8'd147; b = 8'd202;  #10 
a = 8'd147; b = 8'd203;  #10 
a = 8'd147; b = 8'd204;  #10 
a = 8'd147; b = 8'd205;  #10 
a = 8'd147; b = 8'd206;  #10 
a = 8'd147; b = 8'd207;  #10 
a = 8'd147; b = 8'd208;  #10 
a = 8'd147; b = 8'd209;  #10 
a = 8'd147; b = 8'd210;  #10 
a = 8'd147; b = 8'd211;  #10 
a = 8'd147; b = 8'd212;  #10 
a = 8'd147; b = 8'd213;  #10 
a = 8'd147; b = 8'd214;  #10 
a = 8'd147; b = 8'd215;  #10 
a = 8'd147; b = 8'd216;  #10 
a = 8'd147; b = 8'd217;  #10 
a = 8'd147; b = 8'd218;  #10 
a = 8'd147; b = 8'd219;  #10 
a = 8'd147; b = 8'd220;  #10 
a = 8'd147; b = 8'd221;  #10 
a = 8'd147; b = 8'd222;  #10 
a = 8'd147; b = 8'd223;  #10 
a = 8'd147; b = 8'd224;  #10 
a = 8'd147; b = 8'd225;  #10 
a = 8'd147; b = 8'd226;  #10 
a = 8'd147; b = 8'd227;  #10 
a = 8'd147; b = 8'd228;  #10 
a = 8'd147; b = 8'd229;  #10 
a = 8'd147; b = 8'd230;  #10 
a = 8'd147; b = 8'd231;  #10 
a = 8'd147; b = 8'd232;  #10 
a = 8'd147; b = 8'd233;  #10 
a = 8'd147; b = 8'd234;  #10 
a = 8'd147; b = 8'd235;  #10 
a = 8'd147; b = 8'd236;  #10 
a = 8'd147; b = 8'd237;  #10 
a = 8'd147; b = 8'd238;  #10 
a = 8'd147; b = 8'd239;  #10 
a = 8'd147; b = 8'd240;  #10 
a = 8'd147; b = 8'd241;  #10 
a = 8'd147; b = 8'd242;  #10 
a = 8'd147; b = 8'd243;  #10 
a = 8'd147; b = 8'd244;  #10 
a = 8'd147; b = 8'd245;  #10 
a = 8'd147; b = 8'd246;  #10 
a = 8'd147; b = 8'd247;  #10 
a = 8'd147; b = 8'd248;  #10 
a = 8'd147; b = 8'd249;  #10 
a = 8'd147; b = 8'd250;  #10 
a = 8'd147; b = 8'd251;  #10 
a = 8'd147; b = 8'd252;  #10 
a = 8'd147; b = 8'd253;  #10 
a = 8'd147; b = 8'd254;  #10 
a = 8'd147; b = 8'd255;  #10 
a = 8'd148; b = 8'd0;  #10 
a = 8'd148; b = 8'd1;  #10 
a = 8'd148; b = 8'd2;  #10 
a = 8'd148; b = 8'd3;  #10 
a = 8'd148; b = 8'd4;  #10 
a = 8'd148; b = 8'd5;  #10 
a = 8'd148; b = 8'd6;  #10 
a = 8'd148; b = 8'd7;  #10 
a = 8'd148; b = 8'd8;  #10 
a = 8'd148; b = 8'd9;  #10 
a = 8'd148; b = 8'd10;  #10 
a = 8'd148; b = 8'd11;  #10 
a = 8'd148; b = 8'd12;  #10 
a = 8'd148; b = 8'd13;  #10 
a = 8'd148; b = 8'd14;  #10 
a = 8'd148; b = 8'd15;  #10 
a = 8'd148; b = 8'd16;  #10 
a = 8'd148; b = 8'd17;  #10 
a = 8'd148; b = 8'd18;  #10 
a = 8'd148; b = 8'd19;  #10 
a = 8'd148; b = 8'd20;  #10 
a = 8'd148; b = 8'd21;  #10 
a = 8'd148; b = 8'd22;  #10 
a = 8'd148; b = 8'd23;  #10 
a = 8'd148; b = 8'd24;  #10 
a = 8'd148; b = 8'd25;  #10 
a = 8'd148; b = 8'd26;  #10 
a = 8'd148; b = 8'd27;  #10 
a = 8'd148; b = 8'd28;  #10 
a = 8'd148; b = 8'd29;  #10 
a = 8'd148; b = 8'd30;  #10 
a = 8'd148; b = 8'd31;  #10 
a = 8'd148; b = 8'd32;  #10 
a = 8'd148; b = 8'd33;  #10 
a = 8'd148; b = 8'd34;  #10 
a = 8'd148; b = 8'd35;  #10 
a = 8'd148; b = 8'd36;  #10 
a = 8'd148; b = 8'd37;  #10 
a = 8'd148; b = 8'd38;  #10 
a = 8'd148; b = 8'd39;  #10 
a = 8'd148; b = 8'd40;  #10 
a = 8'd148; b = 8'd41;  #10 
a = 8'd148; b = 8'd42;  #10 
a = 8'd148; b = 8'd43;  #10 
a = 8'd148; b = 8'd44;  #10 
a = 8'd148; b = 8'd45;  #10 
a = 8'd148; b = 8'd46;  #10 
a = 8'd148; b = 8'd47;  #10 
a = 8'd148; b = 8'd48;  #10 
a = 8'd148; b = 8'd49;  #10 
a = 8'd148; b = 8'd50;  #10 
a = 8'd148; b = 8'd51;  #10 
a = 8'd148; b = 8'd52;  #10 
a = 8'd148; b = 8'd53;  #10 
a = 8'd148; b = 8'd54;  #10 
a = 8'd148; b = 8'd55;  #10 
a = 8'd148; b = 8'd56;  #10 
a = 8'd148; b = 8'd57;  #10 
a = 8'd148; b = 8'd58;  #10 
a = 8'd148; b = 8'd59;  #10 
a = 8'd148; b = 8'd60;  #10 
a = 8'd148; b = 8'd61;  #10 
a = 8'd148; b = 8'd62;  #10 
a = 8'd148; b = 8'd63;  #10 
a = 8'd148; b = 8'd64;  #10 
a = 8'd148; b = 8'd65;  #10 
a = 8'd148; b = 8'd66;  #10 
a = 8'd148; b = 8'd67;  #10 
a = 8'd148; b = 8'd68;  #10 
a = 8'd148; b = 8'd69;  #10 
a = 8'd148; b = 8'd70;  #10 
a = 8'd148; b = 8'd71;  #10 
a = 8'd148; b = 8'd72;  #10 
a = 8'd148; b = 8'd73;  #10 
a = 8'd148; b = 8'd74;  #10 
a = 8'd148; b = 8'd75;  #10 
a = 8'd148; b = 8'd76;  #10 
a = 8'd148; b = 8'd77;  #10 
a = 8'd148; b = 8'd78;  #10 
a = 8'd148; b = 8'd79;  #10 
a = 8'd148; b = 8'd80;  #10 
a = 8'd148; b = 8'd81;  #10 
a = 8'd148; b = 8'd82;  #10 
a = 8'd148; b = 8'd83;  #10 
a = 8'd148; b = 8'd84;  #10 
a = 8'd148; b = 8'd85;  #10 
a = 8'd148; b = 8'd86;  #10 
a = 8'd148; b = 8'd87;  #10 
a = 8'd148; b = 8'd88;  #10 
a = 8'd148; b = 8'd89;  #10 
a = 8'd148; b = 8'd90;  #10 
a = 8'd148; b = 8'd91;  #10 
a = 8'd148; b = 8'd92;  #10 
a = 8'd148; b = 8'd93;  #10 
a = 8'd148; b = 8'd94;  #10 
a = 8'd148; b = 8'd95;  #10 
a = 8'd148; b = 8'd96;  #10 
a = 8'd148; b = 8'd97;  #10 
a = 8'd148; b = 8'd98;  #10 
a = 8'd148; b = 8'd99;  #10 
a = 8'd148; b = 8'd100;  #10 
a = 8'd148; b = 8'd101;  #10 
a = 8'd148; b = 8'd102;  #10 
a = 8'd148; b = 8'd103;  #10 
a = 8'd148; b = 8'd104;  #10 
a = 8'd148; b = 8'd105;  #10 
a = 8'd148; b = 8'd106;  #10 
a = 8'd148; b = 8'd107;  #10 
a = 8'd148; b = 8'd108;  #10 
a = 8'd148; b = 8'd109;  #10 
a = 8'd148; b = 8'd110;  #10 
a = 8'd148; b = 8'd111;  #10 
a = 8'd148; b = 8'd112;  #10 
a = 8'd148; b = 8'd113;  #10 
a = 8'd148; b = 8'd114;  #10 
a = 8'd148; b = 8'd115;  #10 
a = 8'd148; b = 8'd116;  #10 
a = 8'd148; b = 8'd117;  #10 
a = 8'd148; b = 8'd118;  #10 
a = 8'd148; b = 8'd119;  #10 
a = 8'd148; b = 8'd120;  #10 
a = 8'd148; b = 8'd121;  #10 
a = 8'd148; b = 8'd122;  #10 
a = 8'd148; b = 8'd123;  #10 
a = 8'd148; b = 8'd124;  #10 
a = 8'd148; b = 8'd125;  #10 
a = 8'd148; b = 8'd126;  #10 
a = 8'd148; b = 8'd127;  #10 
a = 8'd148; b = 8'd128;  #10 
a = 8'd148; b = 8'd129;  #10 
a = 8'd148; b = 8'd130;  #10 
a = 8'd148; b = 8'd131;  #10 
a = 8'd148; b = 8'd132;  #10 
a = 8'd148; b = 8'd133;  #10 
a = 8'd148; b = 8'd134;  #10 
a = 8'd148; b = 8'd135;  #10 
a = 8'd148; b = 8'd136;  #10 
a = 8'd148; b = 8'd137;  #10 
a = 8'd148; b = 8'd138;  #10 
a = 8'd148; b = 8'd139;  #10 
a = 8'd148; b = 8'd140;  #10 
a = 8'd148; b = 8'd141;  #10 
a = 8'd148; b = 8'd142;  #10 
a = 8'd148; b = 8'd143;  #10 
a = 8'd148; b = 8'd144;  #10 
a = 8'd148; b = 8'd145;  #10 
a = 8'd148; b = 8'd146;  #10 
a = 8'd148; b = 8'd147;  #10 
a = 8'd148; b = 8'd148;  #10 
a = 8'd148; b = 8'd149;  #10 
a = 8'd148; b = 8'd150;  #10 
a = 8'd148; b = 8'd151;  #10 
a = 8'd148; b = 8'd152;  #10 
a = 8'd148; b = 8'd153;  #10 
a = 8'd148; b = 8'd154;  #10 
a = 8'd148; b = 8'd155;  #10 
a = 8'd148; b = 8'd156;  #10 
a = 8'd148; b = 8'd157;  #10 
a = 8'd148; b = 8'd158;  #10 
a = 8'd148; b = 8'd159;  #10 
a = 8'd148; b = 8'd160;  #10 
a = 8'd148; b = 8'd161;  #10 
a = 8'd148; b = 8'd162;  #10 
a = 8'd148; b = 8'd163;  #10 
a = 8'd148; b = 8'd164;  #10 
a = 8'd148; b = 8'd165;  #10 
a = 8'd148; b = 8'd166;  #10 
a = 8'd148; b = 8'd167;  #10 
a = 8'd148; b = 8'd168;  #10 
a = 8'd148; b = 8'd169;  #10 
a = 8'd148; b = 8'd170;  #10 
a = 8'd148; b = 8'd171;  #10 
a = 8'd148; b = 8'd172;  #10 
a = 8'd148; b = 8'd173;  #10 
a = 8'd148; b = 8'd174;  #10 
a = 8'd148; b = 8'd175;  #10 
a = 8'd148; b = 8'd176;  #10 
a = 8'd148; b = 8'd177;  #10 
a = 8'd148; b = 8'd178;  #10 
a = 8'd148; b = 8'd179;  #10 
a = 8'd148; b = 8'd180;  #10 
a = 8'd148; b = 8'd181;  #10 
a = 8'd148; b = 8'd182;  #10 
a = 8'd148; b = 8'd183;  #10 
a = 8'd148; b = 8'd184;  #10 
a = 8'd148; b = 8'd185;  #10 
a = 8'd148; b = 8'd186;  #10 
a = 8'd148; b = 8'd187;  #10 
a = 8'd148; b = 8'd188;  #10 
a = 8'd148; b = 8'd189;  #10 
a = 8'd148; b = 8'd190;  #10 
a = 8'd148; b = 8'd191;  #10 
a = 8'd148; b = 8'd192;  #10 
a = 8'd148; b = 8'd193;  #10 
a = 8'd148; b = 8'd194;  #10 
a = 8'd148; b = 8'd195;  #10 
a = 8'd148; b = 8'd196;  #10 
a = 8'd148; b = 8'd197;  #10 
a = 8'd148; b = 8'd198;  #10 
a = 8'd148; b = 8'd199;  #10 
a = 8'd148; b = 8'd200;  #10 
a = 8'd148; b = 8'd201;  #10 
a = 8'd148; b = 8'd202;  #10 
a = 8'd148; b = 8'd203;  #10 
a = 8'd148; b = 8'd204;  #10 
a = 8'd148; b = 8'd205;  #10 
a = 8'd148; b = 8'd206;  #10 
a = 8'd148; b = 8'd207;  #10 
a = 8'd148; b = 8'd208;  #10 
a = 8'd148; b = 8'd209;  #10 
a = 8'd148; b = 8'd210;  #10 
a = 8'd148; b = 8'd211;  #10 
a = 8'd148; b = 8'd212;  #10 
a = 8'd148; b = 8'd213;  #10 
a = 8'd148; b = 8'd214;  #10 
a = 8'd148; b = 8'd215;  #10 
a = 8'd148; b = 8'd216;  #10 
a = 8'd148; b = 8'd217;  #10 
a = 8'd148; b = 8'd218;  #10 
a = 8'd148; b = 8'd219;  #10 
a = 8'd148; b = 8'd220;  #10 
a = 8'd148; b = 8'd221;  #10 
a = 8'd148; b = 8'd222;  #10 
a = 8'd148; b = 8'd223;  #10 
a = 8'd148; b = 8'd224;  #10 
a = 8'd148; b = 8'd225;  #10 
a = 8'd148; b = 8'd226;  #10 
a = 8'd148; b = 8'd227;  #10 
a = 8'd148; b = 8'd228;  #10 
a = 8'd148; b = 8'd229;  #10 
a = 8'd148; b = 8'd230;  #10 
a = 8'd148; b = 8'd231;  #10 
a = 8'd148; b = 8'd232;  #10 
a = 8'd148; b = 8'd233;  #10 
a = 8'd148; b = 8'd234;  #10 
a = 8'd148; b = 8'd235;  #10 
a = 8'd148; b = 8'd236;  #10 
a = 8'd148; b = 8'd237;  #10 
a = 8'd148; b = 8'd238;  #10 
a = 8'd148; b = 8'd239;  #10 
a = 8'd148; b = 8'd240;  #10 
a = 8'd148; b = 8'd241;  #10 
a = 8'd148; b = 8'd242;  #10 
a = 8'd148; b = 8'd243;  #10 
a = 8'd148; b = 8'd244;  #10 
a = 8'd148; b = 8'd245;  #10 
a = 8'd148; b = 8'd246;  #10 
a = 8'd148; b = 8'd247;  #10 
a = 8'd148; b = 8'd248;  #10 
a = 8'd148; b = 8'd249;  #10 
a = 8'd148; b = 8'd250;  #10 
a = 8'd148; b = 8'd251;  #10 
a = 8'd148; b = 8'd252;  #10 
a = 8'd148; b = 8'd253;  #10 
a = 8'd148; b = 8'd254;  #10 
a = 8'd148; b = 8'd255;  #10 
a = 8'd149; b = 8'd0;  #10 
a = 8'd149; b = 8'd1;  #10 
a = 8'd149; b = 8'd2;  #10 
a = 8'd149; b = 8'd3;  #10 
a = 8'd149; b = 8'd4;  #10 
a = 8'd149; b = 8'd5;  #10 
a = 8'd149; b = 8'd6;  #10 
a = 8'd149; b = 8'd7;  #10 
a = 8'd149; b = 8'd8;  #10 
a = 8'd149; b = 8'd9;  #10 
a = 8'd149; b = 8'd10;  #10 
a = 8'd149; b = 8'd11;  #10 
a = 8'd149; b = 8'd12;  #10 
a = 8'd149; b = 8'd13;  #10 
a = 8'd149; b = 8'd14;  #10 
a = 8'd149; b = 8'd15;  #10 
a = 8'd149; b = 8'd16;  #10 
a = 8'd149; b = 8'd17;  #10 
a = 8'd149; b = 8'd18;  #10 
a = 8'd149; b = 8'd19;  #10 
a = 8'd149; b = 8'd20;  #10 
a = 8'd149; b = 8'd21;  #10 
a = 8'd149; b = 8'd22;  #10 
a = 8'd149; b = 8'd23;  #10 
a = 8'd149; b = 8'd24;  #10 
a = 8'd149; b = 8'd25;  #10 
a = 8'd149; b = 8'd26;  #10 
a = 8'd149; b = 8'd27;  #10 
a = 8'd149; b = 8'd28;  #10 
a = 8'd149; b = 8'd29;  #10 
a = 8'd149; b = 8'd30;  #10 
a = 8'd149; b = 8'd31;  #10 
a = 8'd149; b = 8'd32;  #10 
a = 8'd149; b = 8'd33;  #10 
a = 8'd149; b = 8'd34;  #10 
a = 8'd149; b = 8'd35;  #10 
a = 8'd149; b = 8'd36;  #10 
a = 8'd149; b = 8'd37;  #10 
a = 8'd149; b = 8'd38;  #10 
a = 8'd149; b = 8'd39;  #10 
a = 8'd149; b = 8'd40;  #10 
a = 8'd149; b = 8'd41;  #10 
a = 8'd149; b = 8'd42;  #10 
a = 8'd149; b = 8'd43;  #10 
a = 8'd149; b = 8'd44;  #10 
a = 8'd149; b = 8'd45;  #10 
a = 8'd149; b = 8'd46;  #10 
a = 8'd149; b = 8'd47;  #10 
a = 8'd149; b = 8'd48;  #10 
a = 8'd149; b = 8'd49;  #10 
a = 8'd149; b = 8'd50;  #10 
a = 8'd149; b = 8'd51;  #10 
a = 8'd149; b = 8'd52;  #10 
a = 8'd149; b = 8'd53;  #10 
a = 8'd149; b = 8'd54;  #10 
a = 8'd149; b = 8'd55;  #10 
a = 8'd149; b = 8'd56;  #10 
a = 8'd149; b = 8'd57;  #10 
a = 8'd149; b = 8'd58;  #10 
a = 8'd149; b = 8'd59;  #10 
a = 8'd149; b = 8'd60;  #10 
a = 8'd149; b = 8'd61;  #10 
a = 8'd149; b = 8'd62;  #10 
a = 8'd149; b = 8'd63;  #10 
a = 8'd149; b = 8'd64;  #10 
a = 8'd149; b = 8'd65;  #10 
a = 8'd149; b = 8'd66;  #10 
a = 8'd149; b = 8'd67;  #10 
a = 8'd149; b = 8'd68;  #10 
a = 8'd149; b = 8'd69;  #10 
a = 8'd149; b = 8'd70;  #10 
a = 8'd149; b = 8'd71;  #10 
a = 8'd149; b = 8'd72;  #10 
a = 8'd149; b = 8'd73;  #10 
a = 8'd149; b = 8'd74;  #10 
a = 8'd149; b = 8'd75;  #10 
a = 8'd149; b = 8'd76;  #10 
a = 8'd149; b = 8'd77;  #10 
a = 8'd149; b = 8'd78;  #10 
a = 8'd149; b = 8'd79;  #10 
a = 8'd149; b = 8'd80;  #10 
a = 8'd149; b = 8'd81;  #10 
a = 8'd149; b = 8'd82;  #10 
a = 8'd149; b = 8'd83;  #10 
a = 8'd149; b = 8'd84;  #10 
a = 8'd149; b = 8'd85;  #10 
a = 8'd149; b = 8'd86;  #10 
a = 8'd149; b = 8'd87;  #10 
a = 8'd149; b = 8'd88;  #10 
a = 8'd149; b = 8'd89;  #10 
a = 8'd149; b = 8'd90;  #10 
a = 8'd149; b = 8'd91;  #10 
a = 8'd149; b = 8'd92;  #10 
a = 8'd149; b = 8'd93;  #10 
a = 8'd149; b = 8'd94;  #10 
a = 8'd149; b = 8'd95;  #10 
a = 8'd149; b = 8'd96;  #10 
a = 8'd149; b = 8'd97;  #10 
a = 8'd149; b = 8'd98;  #10 
a = 8'd149; b = 8'd99;  #10 
a = 8'd149; b = 8'd100;  #10 
a = 8'd149; b = 8'd101;  #10 
a = 8'd149; b = 8'd102;  #10 
a = 8'd149; b = 8'd103;  #10 
a = 8'd149; b = 8'd104;  #10 
a = 8'd149; b = 8'd105;  #10 
a = 8'd149; b = 8'd106;  #10 
a = 8'd149; b = 8'd107;  #10 
a = 8'd149; b = 8'd108;  #10 
a = 8'd149; b = 8'd109;  #10 
a = 8'd149; b = 8'd110;  #10 
a = 8'd149; b = 8'd111;  #10 
a = 8'd149; b = 8'd112;  #10 
a = 8'd149; b = 8'd113;  #10 
a = 8'd149; b = 8'd114;  #10 
a = 8'd149; b = 8'd115;  #10 
a = 8'd149; b = 8'd116;  #10 
a = 8'd149; b = 8'd117;  #10 
a = 8'd149; b = 8'd118;  #10 
a = 8'd149; b = 8'd119;  #10 
a = 8'd149; b = 8'd120;  #10 
a = 8'd149; b = 8'd121;  #10 
a = 8'd149; b = 8'd122;  #10 
a = 8'd149; b = 8'd123;  #10 
a = 8'd149; b = 8'd124;  #10 
a = 8'd149; b = 8'd125;  #10 
a = 8'd149; b = 8'd126;  #10 
a = 8'd149; b = 8'd127;  #10 
a = 8'd149; b = 8'd128;  #10 
a = 8'd149; b = 8'd129;  #10 
a = 8'd149; b = 8'd130;  #10 
a = 8'd149; b = 8'd131;  #10 
a = 8'd149; b = 8'd132;  #10 
a = 8'd149; b = 8'd133;  #10 
a = 8'd149; b = 8'd134;  #10 
a = 8'd149; b = 8'd135;  #10 
a = 8'd149; b = 8'd136;  #10 
a = 8'd149; b = 8'd137;  #10 
a = 8'd149; b = 8'd138;  #10 
a = 8'd149; b = 8'd139;  #10 
a = 8'd149; b = 8'd140;  #10 
a = 8'd149; b = 8'd141;  #10 
a = 8'd149; b = 8'd142;  #10 
a = 8'd149; b = 8'd143;  #10 
a = 8'd149; b = 8'd144;  #10 
a = 8'd149; b = 8'd145;  #10 
a = 8'd149; b = 8'd146;  #10 
a = 8'd149; b = 8'd147;  #10 
a = 8'd149; b = 8'd148;  #10 
a = 8'd149; b = 8'd149;  #10 
a = 8'd149; b = 8'd150;  #10 
a = 8'd149; b = 8'd151;  #10 
a = 8'd149; b = 8'd152;  #10 
a = 8'd149; b = 8'd153;  #10 
a = 8'd149; b = 8'd154;  #10 
a = 8'd149; b = 8'd155;  #10 
a = 8'd149; b = 8'd156;  #10 
a = 8'd149; b = 8'd157;  #10 
a = 8'd149; b = 8'd158;  #10 
a = 8'd149; b = 8'd159;  #10 
a = 8'd149; b = 8'd160;  #10 
a = 8'd149; b = 8'd161;  #10 
a = 8'd149; b = 8'd162;  #10 
a = 8'd149; b = 8'd163;  #10 
a = 8'd149; b = 8'd164;  #10 
a = 8'd149; b = 8'd165;  #10 
a = 8'd149; b = 8'd166;  #10 
a = 8'd149; b = 8'd167;  #10 
a = 8'd149; b = 8'd168;  #10 
a = 8'd149; b = 8'd169;  #10 
a = 8'd149; b = 8'd170;  #10 
a = 8'd149; b = 8'd171;  #10 
a = 8'd149; b = 8'd172;  #10 
a = 8'd149; b = 8'd173;  #10 
a = 8'd149; b = 8'd174;  #10 
a = 8'd149; b = 8'd175;  #10 
a = 8'd149; b = 8'd176;  #10 
a = 8'd149; b = 8'd177;  #10 
a = 8'd149; b = 8'd178;  #10 
a = 8'd149; b = 8'd179;  #10 
a = 8'd149; b = 8'd180;  #10 
a = 8'd149; b = 8'd181;  #10 
a = 8'd149; b = 8'd182;  #10 
a = 8'd149; b = 8'd183;  #10 
a = 8'd149; b = 8'd184;  #10 
a = 8'd149; b = 8'd185;  #10 
a = 8'd149; b = 8'd186;  #10 
a = 8'd149; b = 8'd187;  #10 
a = 8'd149; b = 8'd188;  #10 
a = 8'd149; b = 8'd189;  #10 
a = 8'd149; b = 8'd190;  #10 
a = 8'd149; b = 8'd191;  #10 
a = 8'd149; b = 8'd192;  #10 
a = 8'd149; b = 8'd193;  #10 
a = 8'd149; b = 8'd194;  #10 
a = 8'd149; b = 8'd195;  #10 
a = 8'd149; b = 8'd196;  #10 
a = 8'd149; b = 8'd197;  #10 
a = 8'd149; b = 8'd198;  #10 
a = 8'd149; b = 8'd199;  #10 
a = 8'd149; b = 8'd200;  #10 
a = 8'd149; b = 8'd201;  #10 
a = 8'd149; b = 8'd202;  #10 
a = 8'd149; b = 8'd203;  #10 
a = 8'd149; b = 8'd204;  #10 
a = 8'd149; b = 8'd205;  #10 
a = 8'd149; b = 8'd206;  #10 
a = 8'd149; b = 8'd207;  #10 
a = 8'd149; b = 8'd208;  #10 
a = 8'd149; b = 8'd209;  #10 
a = 8'd149; b = 8'd210;  #10 
a = 8'd149; b = 8'd211;  #10 
a = 8'd149; b = 8'd212;  #10 
a = 8'd149; b = 8'd213;  #10 
a = 8'd149; b = 8'd214;  #10 
a = 8'd149; b = 8'd215;  #10 
a = 8'd149; b = 8'd216;  #10 
a = 8'd149; b = 8'd217;  #10 
a = 8'd149; b = 8'd218;  #10 
a = 8'd149; b = 8'd219;  #10 
a = 8'd149; b = 8'd220;  #10 
a = 8'd149; b = 8'd221;  #10 
a = 8'd149; b = 8'd222;  #10 
a = 8'd149; b = 8'd223;  #10 
a = 8'd149; b = 8'd224;  #10 
a = 8'd149; b = 8'd225;  #10 
a = 8'd149; b = 8'd226;  #10 
a = 8'd149; b = 8'd227;  #10 
a = 8'd149; b = 8'd228;  #10 
a = 8'd149; b = 8'd229;  #10 
a = 8'd149; b = 8'd230;  #10 
a = 8'd149; b = 8'd231;  #10 
a = 8'd149; b = 8'd232;  #10 
a = 8'd149; b = 8'd233;  #10 
a = 8'd149; b = 8'd234;  #10 
a = 8'd149; b = 8'd235;  #10 
a = 8'd149; b = 8'd236;  #10 
a = 8'd149; b = 8'd237;  #10 
a = 8'd149; b = 8'd238;  #10 
a = 8'd149; b = 8'd239;  #10 
a = 8'd149; b = 8'd240;  #10 
a = 8'd149; b = 8'd241;  #10 
a = 8'd149; b = 8'd242;  #10 
a = 8'd149; b = 8'd243;  #10 
a = 8'd149; b = 8'd244;  #10 
a = 8'd149; b = 8'd245;  #10 
a = 8'd149; b = 8'd246;  #10 
a = 8'd149; b = 8'd247;  #10 
a = 8'd149; b = 8'd248;  #10 
a = 8'd149; b = 8'd249;  #10 
a = 8'd149; b = 8'd250;  #10 
a = 8'd149; b = 8'd251;  #10 
a = 8'd149; b = 8'd252;  #10 
a = 8'd149; b = 8'd253;  #10 
a = 8'd149; b = 8'd254;  #10 
a = 8'd149; b = 8'd255;  #10 
a = 8'd150; b = 8'd0;  #10 
a = 8'd150; b = 8'd1;  #10 
a = 8'd150; b = 8'd2;  #10 
a = 8'd150; b = 8'd3;  #10 
a = 8'd150; b = 8'd4;  #10 
a = 8'd150; b = 8'd5;  #10 
a = 8'd150; b = 8'd6;  #10 
a = 8'd150; b = 8'd7;  #10 
a = 8'd150; b = 8'd8;  #10 
a = 8'd150; b = 8'd9;  #10 
a = 8'd150; b = 8'd10;  #10 
a = 8'd150; b = 8'd11;  #10 
a = 8'd150; b = 8'd12;  #10 
a = 8'd150; b = 8'd13;  #10 
a = 8'd150; b = 8'd14;  #10 
a = 8'd150; b = 8'd15;  #10 
a = 8'd150; b = 8'd16;  #10 
a = 8'd150; b = 8'd17;  #10 
a = 8'd150; b = 8'd18;  #10 
a = 8'd150; b = 8'd19;  #10 
a = 8'd150; b = 8'd20;  #10 
a = 8'd150; b = 8'd21;  #10 
a = 8'd150; b = 8'd22;  #10 
a = 8'd150; b = 8'd23;  #10 
a = 8'd150; b = 8'd24;  #10 
a = 8'd150; b = 8'd25;  #10 
a = 8'd150; b = 8'd26;  #10 
a = 8'd150; b = 8'd27;  #10 
a = 8'd150; b = 8'd28;  #10 
a = 8'd150; b = 8'd29;  #10 
a = 8'd150; b = 8'd30;  #10 
a = 8'd150; b = 8'd31;  #10 
a = 8'd150; b = 8'd32;  #10 
a = 8'd150; b = 8'd33;  #10 
a = 8'd150; b = 8'd34;  #10 
a = 8'd150; b = 8'd35;  #10 
a = 8'd150; b = 8'd36;  #10 
a = 8'd150; b = 8'd37;  #10 
a = 8'd150; b = 8'd38;  #10 
a = 8'd150; b = 8'd39;  #10 
a = 8'd150; b = 8'd40;  #10 
a = 8'd150; b = 8'd41;  #10 
a = 8'd150; b = 8'd42;  #10 
a = 8'd150; b = 8'd43;  #10 
a = 8'd150; b = 8'd44;  #10 
a = 8'd150; b = 8'd45;  #10 
a = 8'd150; b = 8'd46;  #10 
a = 8'd150; b = 8'd47;  #10 
a = 8'd150; b = 8'd48;  #10 
a = 8'd150; b = 8'd49;  #10 
a = 8'd150; b = 8'd50;  #10 
a = 8'd150; b = 8'd51;  #10 
a = 8'd150; b = 8'd52;  #10 
a = 8'd150; b = 8'd53;  #10 
a = 8'd150; b = 8'd54;  #10 
a = 8'd150; b = 8'd55;  #10 
a = 8'd150; b = 8'd56;  #10 
a = 8'd150; b = 8'd57;  #10 
a = 8'd150; b = 8'd58;  #10 
a = 8'd150; b = 8'd59;  #10 
a = 8'd150; b = 8'd60;  #10 
a = 8'd150; b = 8'd61;  #10 
a = 8'd150; b = 8'd62;  #10 
a = 8'd150; b = 8'd63;  #10 
a = 8'd150; b = 8'd64;  #10 
a = 8'd150; b = 8'd65;  #10 
a = 8'd150; b = 8'd66;  #10 
a = 8'd150; b = 8'd67;  #10 
a = 8'd150; b = 8'd68;  #10 
a = 8'd150; b = 8'd69;  #10 
a = 8'd150; b = 8'd70;  #10 
a = 8'd150; b = 8'd71;  #10 
a = 8'd150; b = 8'd72;  #10 
a = 8'd150; b = 8'd73;  #10 
a = 8'd150; b = 8'd74;  #10 
a = 8'd150; b = 8'd75;  #10 
a = 8'd150; b = 8'd76;  #10 
a = 8'd150; b = 8'd77;  #10 
a = 8'd150; b = 8'd78;  #10 
a = 8'd150; b = 8'd79;  #10 
a = 8'd150; b = 8'd80;  #10 
a = 8'd150; b = 8'd81;  #10 
a = 8'd150; b = 8'd82;  #10 
a = 8'd150; b = 8'd83;  #10 
a = 8'd150; b = 8'd84;  #10 
a = 8'd150; b = 8'd85;  #10 
a = 8'd150; b = 8'd86;  #10 
a = 8'd150; b = 8'd87;  #10 
a = 8'd150; b = 8'd88;  #10 
a = 8'd150; b = 8'd89;  #10 
a = 8'd150; b = 8'd90;  #10 
a = 8'd150; b = 8'd91;  #10 
a = 8'd150; b = 8'd92;  #10 
a = 8'd150; b = 8'd93;  #10 
a = 8'd150; b = 8'd94;  #10 
a = 8'd150; b = 8'd95;  #10 
a = 8'd150; b = 8'd96;  #10 
a = 8'd150; b = 8'd97;  #10 
a = 8'd150; b = 8'd98;  #10 
a = 8'd150; b = 8'd99;  #10 
a = 8'd150; b = 8'd100;  #10 
a = 8'd150; b = 8'd101;  #10 
a = 8'd150; b = 8'd102;  #10 
a = 8'd150; b = 8'd103;  #10 
a = 8'd150; b = 8'd104;  #10 
a = 8'd150; b = 8'd105;  #10 
a = 8'd150; b = 8'd106;  #10 
a = 8'd150; b = 8'd107;  #10 
a = 8'd150; b = 8'd108;  #10 
a = 8'd150; b = 8'd109;  #10 
a = 8'd150; b = 8'd110;  #10 
a = 8'd150; b = 8'd111;  #10 
a = 8'd150; b = 8'd112;  #10 
a = 8'd150; b = 8'd113;  #10 
a = 8'd150; b = 8'd114;  #10 
a = 8'd150; b = 8'd115;  #10 
a = 8'd150; b = 8'd116;  #10 
a = 8'd150; b = 8'd117;  #10 
a = 8'd150; b = 8'd118;  #10 
a = 8'd150; b = 8'd119;  #10 
a = 8'd150; b = 8'd120;  #10 
a = 8'd150; b = 8'd121;  #10 
a = 8'd150; b = 8'd122;  #10 
a = 8'd150; b = 8'd123;  #10 
a = 8'd150; b = 8'd124;  #10 
a = 8'd150; b = 8'd125;  #10 
a = 8'd150; b = 8'd126;  #10 
a = 8'd150; b = 8'd127;  #10 
a = 8'd150; b = 8'd128;  #10 
a = 8'd150; b = 8'd129;  #10 
a = 8'd150; b = 8'd130;  #10 
a = 8'd150; b = 8'd131;  #10 
a = 8'd150; b = 8'd132;  #10 
a = 8'd150; b = 8'd133;  #10 
a = 8'd150; b = 8'd134;  #10 
a = 8'd150; b = 8'd135;  #10 
a = 8'd150; b = 8'd136;  #10 
a = 8'd150; b = 8'd137;  #10 
a = 8'd150; b = 8'd138;  #10 
a = 8'd150; b = 8'd139;  #10 
a = 8'd150; b = 8'd140;  #10 
a = 8'd150; b = 8'd141;  #10 
a = 8'd150; b = 8'd142;  #10 
a = 8'd150; b = 8'd143;  #10 
a = 8'd150; b = 8'd144;  #10 
a = 8'd150; b = 8'd145;  #10 
a = 8'd150; b = 8'd146;  #10 
a = 8'd150; b = 8'd147;  #10 
a = 8'd150; b = 8'd148;  #10 
a = 8'd150; b = 8'd149;  #10 
a = 8'd150; b = 8'd150;  #10 
a = 8'd150; b = 8'd151;  #10 
a = 8'd150; b = 8'd152;  #10 
a = 8'd150; b = 8'd153;  #10 
a = 8'd150; b = 8'd154;  #10 
a = 8'd150; b = 8'd155;  #10 
a = 8'd150; b = 8'd156;  #10 
a = 8'd150; b = 8'd157;  #10 
a = 8'd150; b = 8'd158;  #10 
a = 8'd150; b = 8'd159;  #10 
a = 8'd150; b = 8'd160;  #10 
a = 8'd150; b = 8'd161;  #10 
a = 8'd150; b = 8'd162;  #10 
a = 8'd150; b = 8'd163;  #10 
a = 8'd150; b = 8'd164;  #10 
a = 8'd150; b = 8'd165;  #10 
a = 8'd150; b = 8'd166;  #10 
a = 8'd150; b = 8'd167;  #10 
a = 8'd150; b = 8'd168;  #10 
a = 8'd150; b = 8'd169;  #10 
a = 8'd150; b = 8'd170;  #10 
a = 8'd150; b = 8'd171;  #10 
a = 8'd150; b = 8'd172;  #10 
a = 8'd150; b = 8'd173;  #10 
a = 8'd150; b = 8'd174;  #10 
a = 8'd150; b = 8'd175;  #10 
a = 8'd150; b = 8'd176;  #10 
a = 8'd150; b = 8'd177;  #10 
a = 8'd150; b = 8'd178;  #10 
a = 8'd150; b = 8'd179;  #10 
a = 8'd150; b = 8'd180;  #10 
a = 8'd150; b = 8'd181;  #10 
a = 8'd150; b = 8'd182;  #10 
a = 8'd150; b = 8'd183;  #10 
a = 8'd150; b = 8'd184;  #10 
a = 8'd150; b = 8'd185;  #10 
a = 8'd150; b = 8'd186;  #10 
a = 8'd150; b = 8'd187;  #10 
a = 8'd150; b = 8'd188;  #10 
a = 8'd150; b = 8'd189;  #10 
a = 8'd150; b = 8'd190;  #10 
a = 8'd150; b = 8'd191;  #10 
a = 8'd150; b = 8'd192;  #10 
a = 8'd150; b = 8'd193;  #10 
a = 8'd150; b = 8'd194;  #10 
a = 8'd150; b = 8'd195;  #10 
a = 8'd150; b = 8'd196;  #10 
a = 8'd150; b = 8'd197;  #10 
a = 8'd150; b = 8'd198;  #10 
a = 8'd150; b = 8'd199;  #10 
a = 8'd150; b = 8'd200;  #10 
a = 8'd150; b = 8'd201;  #10 
a = 8'd150; b = 8'd202;  #10 
a = 8'd150; b = 8'd203;  #10 
a = 8'd150; b = 8'd204;  #10 
a = 8'd150; b = 8'd205;  #10 
a = 8'd150; b = 8'd206;  #10 
a = 8'd150; b = 8'd207;  #10 
a = 8'd150; b = 8'd208;  #10 
a = 8'd150; b = 8'd209;  #10 
a = 8'd150; b = 8'd210;  #10 
a = 8'd150; b = 8'd211;  #10 
a = 8'd150; b = 8'd212;  #10 
a = 8'd150; b = 8'd213;  #10 
a = 8'd150; b = 8'd214;  #10 
a = 8'd150; b = 8'd215;  #10 
a = 8'd150; b = 8'd216;  #10 
a = 8'd150; b = 8'd217;  #10 
a = 8'd150; b = 8'd218;  #10 
a = 8'd150; b = 8'd219;  #10 
a = 8'd150; b = 8'd220;  #10 
a = 8'd150; b = 8'd221;  #10 
a = 8'd150; b = 8'd222;  #10 
a = 8'd150; b = 8'd223;  #10 
a = 8'd150; b = 8'd224;  #10 
a = 8'd150; b = 8'd225;  #10 
a = 8'd150; b = 8'd226;  #10 
a = 8'd150; b = 8'd227;  #10 
a = 8'd150; b = 8'd228;  #10 
a = 8'd150; b = 8'd229;  #10 
a = 8'd150; b = 8'd230;  #10 
a = 8'd150; b = 8'd231;  #10 
a = 8'd150; b = 8'd232;  #10 
a = 8'd150; b = 8'd233;  #10 
a = 8'd150; b = 8'd234;  #10 
a = 8'd150; b = 8'd235;  #10 
a = 8'd150; b = 8'd236;  #10 
a = 8'd150; b = 8'd237;  #10 
a = 8'd150; b = 8'd238;  #10 
a = 8'd150; b = 8'd239;  #10 
a = 8'd150; b = 8'd240;  #10 
a = 8'd150; b = 8'd241;  #10 
a = 8'd150; b = 8'd242;  #10 
a = 8'd150; b = 8'd243;  #10 
a = 8'd150; b = 8'd244;  #10 
a = 8'd150; b = 8'd245;  #10 
a = 8'd150; b = 8'd246;  #10 
a = 8'd150; b = 8'd247;  #10 
a = 8'd150; b = 8'd248;  #10 
a = 8'd150; b = 8'd249;  #10 
a = 8'd150; b = 8'd250;  #10 
a = 8'd150; b = 8'd251;  #10 
a = 8'd150; b = 8'd252;  #10 
a = 8'd150; b = 8'd253;  #10 
a = 8'd150; b = 8'd254;  #10 
a = 8'd150; b = 8'd255;  #10 
a = 8'd151; b = 8'd0;  #10 
a = 8'd151; b = 8'd1;  #10 
a = 8'd151; b = 8'd2;  #10 
a = 8'd151; b = 8'd3;  #10 
a = 8'd151; b = 8'd4;  #10 
a = 8'd151; b = 8'd5;  #10 
a = 8'd151; b = 8'd6;  #10 
a = 8'd151; b = 8'd7;  #10 
a = 8'd151; b = 8'd8;  #10 
a = 8'd151; b = 8'd9;  #10 
a = 8'd151; b = 8'd10;  #10 
a = 8'd151; b = 8'd11;  #10 
a = 8'd151; b = 8'd12;  #10 
a = 8'd151; b = 8'd13;  #10 
a = 8'd151; b = 8'd14;  #10 
a = 8'd151; b = 8'd15;  #10 
a = 8'd151; b = 8'd16;  #10 
a = 8'd151; b = 8'd17;  #10 
a = 8'd151; b = 8'd18;  #10 
a = 8'd151; b = 8'd19;  #10 
a = 8'd151; b = 8'd20;  #10 
a = 8'd151; b = 8'd21;  #10 
a = 8'd151; b = 8'd22;  #10 
a = 8'd151; b = 8'd23;  #10 
a = 8'd151; b = 8'd24;  #10 
a = 8'd151; b = 8'd25;  #10 
a = 8'd151; b = 8'd26;  #10 
a = 8'd151; b = 8'd27;  #10 
a = 8'd151; b = 8'd28;  #10 
a = 8'd151; b = 8'd29;  #10 
a = 8'd151; b = 8'd30;  #10 
a = 8'd151; b = 8'd31;  #10 
a = 8'd151; b = 8'd32;  #10 
a = 8'd151; b = 8'd33;  #10 
a = 8'd151; b = 8'd34;  #10 
a = 8'd151; b = 8'd35;  #10 
a = 8'd151; b = 8'd36;  #10 
a = 8'd151; b = 8'd37;  #10 
a = 8'd151; b = 8'd38;  #10 
a = 8'd151; b = 8'd39;  #10 
a = 8'd151; b = 8'd40;  #10 
a = 8'd151; b = 8'd41;  #10 
a = 8'd151; b = 8'd42;  #10 
a = 8'd151; b = 8'd43;  #10 
a = 8'd151; b = 8'd44;  #10 
a = 8'd151; b = 8'd45;  #10 
a = 8'd151; b = 8'd46;  #10 
a = 8'd151; b = 8'd47;  #10 
a = 8'd151; b = 8'd48;  #10 
a = 8'd151; b = 8'd49;  #10 
a = 8'd151; b = 8'd50;  #10 
a = 8'd151; b = 8'd51;  #10 
a = 8'd151; b = 8'd52;  #10 
a = 8'd151; b = 8'd53;  #10 
a = 8'd151; b = 8'd54;  #10 
a = 8'd151; b = 8'd55;  #10 
a = 8'd151; b = 8'd56;  #10 
a = 8'd151; b = 8'd57;  #10 
a = 8'd151; b = 8'd58;  #10 
a = 8'd151; b = 8'd59;  #10 
a = 8'd151; b = 8'd60;  #10 
a = 8'd151; b = 8'd61;  #10 
a = 8'd151; b = 8'd62;  #10 
a = 8'd151; b = 8'd63;  #10 
a = 8'd151; b = 8'd64;  #10 
a = 8'd151; b = 8'd65;  #10 
a = 8'd151; b = 8'd66;  #10 
a = 8'd151; b = 8'd67;  #10 
a = 8'd151; b = 8'd68;  #10 
a = 8'd151; b = 8'd69;  #10 
a = 8'd151; b = 8'd70;  #10 
a = 8'd151; b = 8'd71;  #10 
a = 8'd151; b = 8'd72;  #10 
a = 8'd151; b = 8'd73;  #10 
a = 8'd151; b = 8'd74;  #10 
a = 8'd151; b = 8'd75;  #10 
a = 8'd151; b = 8'd76;  #10 
a = 8'd151; b = 8'd77;  #10 
a = 8'd151; b = 8'd78;  #10 
a = 8'd151; b = 8'd79;  #10 
a = 8'd151; b = 8'd80;  #10 
a = 8'd151; b = 8'd81;  #10 
a = 8'd151; b = 8'd82;  #10 
a = 8'd151; b = 8'd83;  #10 
a = 8'd151; b = 8'd84;  #10 
a = 8'd151; b = 8'd85;  #10 
a = 8'd151; b = 8'd86;  #10 
a = 8'd151; b = 8'd87;  #10 
a = 8'd151; b = 8'd88;  #10 
a = 8'd151; b = 8'd89;  #10 
a = 8'd151; b = 8'd90;  #10 
a = 8'd151; b = 8'd91;  #10 
a = 8'd151; b = 8'd92;  #10 
a = 8'd151; b = 8'd93;  #10 
a = 8'd151; b = 8'd94;  #10 
a = 8'd151; b = 8'd95;  #10 
a = 8'd151; b = 8'd96;  #10 
a = 8'd151; b = 8'd97;  #10 
a = 8'd151; b = 8'd98;  #10 
a = 8'd151; b = 8'd99;  #10 
a = 8'd151; b = 8'd100;  #10 
a = 8'd151; b = 8'd101;  #10 
a = 8'd151; b = 8'd102;  #10 
a = 8'd151; b = 8'd103;  #10 
a = 8'd151; b = 8'd104;  #10 
a = 8'd151; b = 8'd105;  #10 
a = 8'd151; b = 8'd106;  #10 
a = 8'd151; b = 8'd107;  #10 
a = 8'd151; b = 8'd108;  #10 
a = 8'd151; b = 8'd109;  #10 
a = 8'd151; b = 8'd110;  #10 
a = 8'd151; b = 8'd111;  #10 
a = 8'd151; b = 8'd112;  #10 
a = 8'd151; b = 8'd113;  #10 
a = 8'd151; b = 8'd114;  #10 
a = 8'd151; b = 8'd115;  #10 
a = 8'd151; b = 8'd116;  #10 
a = 8'd151; b = 8'd117;  #10 
a = 8'd151; b = 8'd118;  #10 
a = 8'd151; b = 8'd119;  #10 
a = 8'd151; b = 8'd120;  #10 
a = 8'd151; b = 8'd121;  #10 
a = 8'd151; b = 8'd122;  #10 
a = 8'd151; b = 8'd123;  #10 
a = 8'd151; b = 8'd124;  #10 
a = 8'd151; b = 8'd125;  #10 
a = 8'd151; b = 8'd126;  #10 
a = 8'd151; b = 8'd127;  #10 
a = 8'd151; b = 8'd128;  #10 
a = 8'd151; b = 8'd129;  #10 
a = 8'd151; b = 8'd130;  #10 
a = 8'd151; b = 8'd131;  #10 
a = 8'd151; b = 8'd132;  #10 
a = 8'd151; b = 8'd133;  #10 
a = 8'd151; b = 8'd134;  #10 
a = 8'd151; b = 8'd135;  #10 
a = 8'd151; b = 8'd136;  #10 
a = 8'd151; b = 8'd137;  #10 
a = 8'd151; b = 8'd138;  #10 
a = 8'd151; b = 8'd139;  #10 
a = 8'd151; b = 8'd140;  #10 
a = 8'd151; b = 8'd141;  #10 
a = 8'd151; b = 8'd142;  #10 
a = 8'd151; b = 8'd143;  #10 
a = 8'd151; b = 8'd144;  #10 
a = 8'd151; b = 8'd145;  #10 
a = 8'd151; b = 8'd146;  #10 
a = 8'd151; b = 8'd147;  #10 
a = 8'd151; b = 8'd148;  #10 
a = 8'd151; b = 8'd149;  #10 
a = 8'd151; b = 8'd150;  #10 
a = 8'd151; b = 8'd151;  #10 
a = 8'd151; b = 8'd152;  #10 
a = 8'd151; b = 8'd153;  #10 
a = 8'd151; b = 8'd154;  #10 
a = 8'd151; b = 8'd155;  #10 
a = 8'd151; b = 8'd156;  #10 
a = 8'd151; b = 8'd157;  #10 
a = 8'd151; b = 8'd158;  #10 
a = 8'd151; b = 8'd159;  #10 
a = 8'd151; b = 8'd160;  #10 
a = 8'd151; b = 8'd161;  #10 
a = 8'd151; b = 8'd162;  #10 
a = 8'd151; b = 8'd163;  #10 
a = 8'd151; b = 8'd164;  #10 
a = 8'd151; b = 8'd165;  #10 
a = 8'd151; b = 8'd166;  #10 
a = 8'd151; b = 8'd167;  #10 
a = 8'd151; b = 8'd168;  #10 
a = 8'd151; b = 8'd169;  #10 
a = 8'd151; b = 8'd170;  #10 
a = 8'd151; b = 8'd171;  #10 
a = 8'd151; b = 8'd172;  #10 
a = 8'd151; b = 8'd173;  #10 
a = 8'd151; b = 8'd174;  #10 
a = 8'd151; b = 8'd175;  #10 
a = 8'd151; b = 8'd176;  #10 
a = 8'd151; b = 8'd177;  #10 
a = 8'd151; b = 8'd178;  #10 
a = 8'd151; b = 8'd179;  #10 
a = 8'd151; b = 8'd180;  #10 
a = 8'd151; b = 8'd181;  #10 
a = 8'd151; b = 8'd182;  #10 
a = 8'd151; b = 8'd183;  #10 
a = 8'd151; b = 8'd184;  #10 
a = 8'd151; b = 8'd185;  #10 
a = 8'd151; b = 8'd186;  #10 
a = 8'd151; b = 8'd187;  #10 
a = 8'd151; b = 8'd188;  #10 
a = 8'd151; b = 8'd189;  #10 
a = 8'd151; b = 8'd190;  #10 
a = 8'd151; b = 8'd191;  #10 
a = 8'd151; b = 8'd192;  #10 
a = 8'd151; b = 8'd193;  #10 
a = 8'd151; b = 8'd194;  #10 
a = 8'd151; b = 8'd195;  #10 
a = 8'd151; b = 8'd196;  #10 
a = 8'd151; b = 8'd197;  #10 
a = 8'd151; b = 8'd198;  #10 
a = 8'd151; b = 8'd199;  #10 
a = 8'd151; b = 8'd200;  #10 
a = 8'd151; b = 8'd201;  #10 
a = 8'd151; b = 8'd202;  #10 
a = 8'd151; b = 8'd203;  #10 
a = 8'd151; b = 8'd204;  #10 
a = 8'd151; b = 8'd205;  #10 
a = 8'd151; b = 8'd206;  #10 
a = 8'd151; b = 8'd207;  #10 
a = 8'd151; b = 8'd208;  #10 
a = 8'd151; b = 8'd209;  #10 
a = 8'd151; b = 8'd210;  #10 
a = 8'd151; b = 8'd211;  #10 
a = 8'd151; b = 8'd212;  #10 
a = 8'd151; b = 8'd213;  #10 
a = 8'd151; b = 8'd214;  #10 
a = 8'd151; b = 8'd215;  #10 
a = 8'd151; b = 8'd216;  #10 
a = 8'd151; b = 8'd217;  #10 
a = 8'd151; b = 8'd218;  #10 
a = 8'd151; b = 8'd219;  #10 
a = 8'd151; b = 8'd220;  #10 
a = 8'd151; b = 8'd221;  #10 
a = 8'd151; b = 8'd222;  #10 
a = 8'd151; b = 8'd223;  #10 
a = 8'd151; b = 8'd224;  #10 
a = 8'd151; b = 8'd225;  #10 
a = 8'd151; b = 8'd226;  #10 
a = 8'd151; b = 8'd227;  #10 
a = 8'd151; b = 8'd228;  #10 
a = 8'd151; b = 8'd229;  #10 
a = 8'd151; b = 8'd230;  #10 
a = 8'd151; b = 8'd231;  #10 
a = 8'd151; b = 8'd232;  #10 
a = 8'd151; b = 8'd233;  #10 
a = 8'd151; b = 8'd234;  #10 
a = 8'd151; b = 8'd235;  #10 
a = 8'd151; b = 8'd236;  #10 
a = 8'd151; b = 8'd237;  #10 
a = 8'd151; b = 8'd238;  #10 
a = 8'd151; b = 8'd239;  #10 
a = 8'd151; b = 8'd240;  #10 
a = 8'd151; b = 8'd241;  #10 
a = 8'd151; b = 8'd242;  #10 
a = 8'd151; b = 8'd243;  #10 
a = 8'd151; b = 8'd244;  #10 
a = 8'd151; b = 8'd245;  #10 
a = 8'd151; b = 8'd246;  #10 
a = 8'd151; b = 8'd247;  #10 
a = 8'd151; b = 8'd248;  #10 
a = 8'd151; b = 8'd249;  #10 
a = 8'd151; b = 8'd250;  #10 
a = 8'd151; b = 8'd251;  #10 
a = 8'd151; b = 8'd252;  #10 
a = 8'd151; b = 8'd253;  #10 
a = 8'd151; b = 8'd254;  #10 
a = 8'd151; b = 8'd255;  #10 
a = 8'd152; b = 8'd0;  #10 
a = 8'd152; b = 8'd1;  #10 
a = 8'd152; b = 8'd2;  #10 
a = 8'd152; b = 8'd3;  #10 
a = 8'd152; b = 8'd4;  #10 
a = 8'd152; b = 8'd5;  #10 
a = 8'd152; b = 8'd6;  #10 
a = 8'd152; b = 8'd7;  #10 
a = 8'd152; b = 8'd8;  #10 
a = 8'd152; b = 8'd9;  #10 
a = 8'd152; b = 8'd10;  #10 
a = 8'd152; b = 8'd11;  #10 
a = 8'd152; b = 8'd12;  #10 
a = 8'd152; b = 8'd13;  #10 
a = 8'd152; b = 8'd14;  #10 
a = 8'd152; b = 8'd15;  #10 
a = 8'd152; b = 8'd16;  #10 
a = 8'd152; b = 8'd17;  #10 
a = 8'd152; b = 8'd18;  #10 
a = 8'd152; b = 8'd19;  #10 
a = 8'd152; b = 8'd20;  #10 
a = 8'd152; b = 8'd21;  #10 
a = 8'd152; b = 8'd22;  #10 
a = 8'd152; b = 8'd23;  #10 
a = 8'd152; b = 8'd24;  #10 
a = 8'd152; b = 8'd25;  #10 
a = 8'd152; b = 8'd26;  #10 
a = 8'd152; b = 8'd27;  #10 
a = 8'd152; b = 8'd28;  #10 
a = 8'd152; b = 8'd29;  #10 
a = 8'd152; b = 8'd30;  #10 
a = 8'd152; b = 8'd31;  #10 
a = 8'd152; b = 8'd32;  #10 
a = 8'd152; b = 8'd33;  #10 
a = 8'd152; b = 8'd34;  #10 
a = 8'd152; b = 8'd35;  #10 
a = 8'd152; b = 8'd36;  #10 
a = 8'd152; b = 8'd37;  #10 
a = 8'd152; b = 8'd38;  #10 
a = 8'd152; b = 8'd39;  #10 
a = 8'd152; b = 8'd40;  #10 
a = 8'd152; b = 8'd41;  #10 
a = 8'd152; b = 8'd42;  #10 
a = 8'd152; b = 8'd43;  #10 
a = 8'd152; b = 8'd44;  #10 
a = 8'd152; b = 8'd45;  #10 
a = 8'd152; b = 8'd46;  #10 
a = 8'd152; b = 8'd47;  #10 
a = 8'd152; b = 8'd48;  #10 
a = 8'd152; b = 8'd49;  #10 
a = 8'd152; b = 8'd50;  #10 
a = 8'd152; b = 8'd51;  #10 
a = 8'd152; b = 8'd52;  #10 
a = 8'd152; b = 8'd53;  #10 
a = 8'd152; b = 8'd54;  #10 
a = 8'd152; b = 8'd55;  #10 
a = 8'd152; b = 8'd56;  #10 
a = 8'd152; b = 8'd57;  #10 
a = 8'd152; b = 8'd58;  #10 
a = 8'd152; b = 8'd59;  #10 
a = 8'd152; b = 8'd60;  #10 
a = 8'd152; b = 8'd61;  #10 
a = 8'd152; b = 8'd62;  #10 
a = 8'd152; b = 8'd63;  #10 
a = 8'd152; b = 8'd64;  #10 
a = 8'd152; b = 8'd65;  #10 
a = 8'd152; b = 8'd66;  #10 
a = 8'd152; b = 8'd67;  #10 
a = 8'd152; b = 8'd68;  #10 
a = 8'd152; b = 8'd69;  #10 
a = 8'd152; b = 8'd70;  #10 
a = 8'd152; b = 8'd71;  #10 
a = 8'd152; b = 8'd72;  #10 
a = 8'd152; b = 8'd73;  #10 
a = 8'd152; b = 8'd74;  #10 
a = 8'd152; b = 8'd75;  #10 
a = 8'd152; b = 8'd76;  #10 
a = 8'd152; b = 8'd77;  #10 
a = 8'd152; b = 8'd78;  #10 
a = 8'd152; b = 8'd79;  #10 
a = 8'd152; b = 8'd80;  #10 
a = 8'd152; b = 8'd81;  #10 
a = 8'd152; b = 8'd82;  #10 
a = 8'd152; b = 8'd83;  #10 
a = 8'd152; b = 8'd84;  #10 
a = 8'd152; b = 8'd85;  #10 
a = 8'd152; b = 8'd86;  #10 
a = 8'd152; b = 8'd87;  #10 
a = 8'd152; b = 8'd88;  #10 
a = 8'd152; b = 8'd89;  #10 
a = 8'd152; b = 8'd90;  #10 
a = 8'd152; b = 8'd91;  #10 
a = 8'd152; b = 8'd92;  #10 
a = 8'd152; b = 8'd93;  #10 
a = 8'd152; b = 8'd94;  #10 
a = 8'd152; b = 8'd95;  #10 
a = 8'd152; b = 8'd96;  #10 
a = 8'd152; b = 8'd97;  #10 
a = 8'd152; b = 8'd98;  #10 
a = 8'd152; b = 8'd99;  #10 
a = 8'd152; b = 8'd100;  #10 
a = 8'd152; b = 8'd101;  #10 
a = 8'd152; b = 8'd102;  #10 
a = 8'd152; b = 8'd103;  #10 
a = 8'd152; b = 8'd104;  #10 
a = 8'd152; b = 8'd105;  #10 
a = 8'd152; b = 8'd106;  #10 
a = 8'd152; b = 8'd107;  #10 
a = 8'd152; b = 8'd108;  #10 
a = 8'd152; b = 8'd109;  #10 
a = 8'd152; b = 8'd110;  #10 
a = 8'd152; b = 8'd111;  #10 
a = 8'd152; b = 8'd112;  #10 
a = 8'd152; b = 8'd113;  #10 
a = 8'd152; b = 8'd114;  #10 
a = 8'd152; b = 8'd115;  #10 
a = 8'd152; b = 8'd116;  #10 
a = 8'd152; b = 8'd117;  #10 
a = 8'd152; b = 8'd118;  #10 
a = 8'd152; b = 8'd119;  #10 
a = 8'd152; b = 8'd120;  #10 
a = 8'd152; b = 8'd121;  #10 
a = 8'd152; b = 8'd122;  #10 
a = 8'd152; b = 8'd123;  #10 
a = 8'd152; b = 8'd124;  #10 
a = 8'd152; b = 8'd125;  #10 
a = 8'd152; b = 8'd126;  #10 
a = 8'd152; b = 8'd127;  #10 
a = 8'd152; b = 8'd128;  #10 
a = 8'd152; b = 8'd129;  #10 
a = 8'd152; b = 8'd130;  #10 
a = 8'd152; b = 8'd131;  #10 
a = 8'd152; b = 8'd132;  #10 
a = 8'd152; b = 8'd133;  #10 
a = 8'd152; b = 8'd134;  #10 
a = 8'd152; b = 8'd135;  #10 
a = 8'd152; b = 8'd136;  #10 
a = 8'd152; b = 8'd137;  #10 
a = 8'd152; b = 8'd138;  #10 
a = 8'd152; b = 8'd139;  #10 
a = 8'd152; b = 8'd140;  #10 
a = 8'd152; b = 8'd141;  #10 
a = 8'd152; b = 8'd142;  #10 
a = 8'd152; b = 8'd143;  #10 
a = 8'd152; b = 8'd144;  #10 
a = 8'd152; b = 8'd145;  #10 
a = 8'd152; b = 8'd146;  #10 
a = 8'd152; b = 8'd147;  #10 
a = 8'd152; b = 8'd148;  #10 
a = 8'd152; b = 8'd149;  #10 
a = 8'd152; b = 8'd150;  #10 
a = 8'd152; b = 8'd151;  #10 
a = 8'd152; b = 8'd152;  #10 
a = 8'd152; b = 8'd153;  #10 
a = 8'd152; b = 8'd154;  #10 
a = 8'd152; b = 8'd155;  #10 
a = 8'd152; b = 8'd156;  #10 
a = 8'd152; b = 8'd157;  #10 
a = 8'd152; b = 8'd158;  #10 
a = 8'd152; b = 8'd159;  #10 
a = 8'd152; b = 8'd160;  #10 
a = 8'd152; b = 8'd161;  #10 
a = 8'd152; b = 8'd162;  #10 
a = 8'd152; b = 8'd163;  #10 
a = 8'd152; b = 8'd164;  #10 
a = 8'd152; b = 8'd165;  #10 
a = 8'd152; b = 8'd166;  #10 
a = 8'd152; b = 8'd167;  #10 
a = 8'd152; b = 8'd168;  #10 
a = 8'd152; b = 8'd169;  #10 
a = 8'd152; b = 8'd170;  #10 
a = 8'd152; b = 8'd171;  #10 
a = 8'd152; b = 8'd172;  #10 
a = 8'd152; b = 8'd173;  #10 
a = 8'd152; b = 8'd174;  #10 
a = 8'd152; b = 8'd175;  #10 
a = 8'd152; b = 8'd176;  #10 
a = 8'd152; b = 8'd177;  #10 
a = 8'd152; b = 8'd178;  #10 
a = 8'd152; b = 8'd179;  #10 
a = 8'd152; b = 8'd180;  #10 
a = 8'd152; b = 8'd181;  #10 
a = 8'd152; b = 8'd182;  #10 
a = 8'd152; b = 8'd183;  #10 
a = 8'd152; b = 8'd184;  #10 
a = 8'd152; b = 8'd185;  #10 
a = 8'd152; b = 8'd186;  #10 
a = 8'd152; b = 8'd187;  #10 
a = 8'd152; b = 8'd188;  #10 
a = 8'd152; b = 8'd189;  #10 
a = 8'd152; b = 8'd190;  #10 
a = 8'd152; b = 8'd191;  #10 
a = 8'd152; b = 8'd192;  #10 
a = 8'd152; b = 8'd193;  #10 
a = 8'd152; b = 8'd194;  #10 
a = 8'd152; b = 8'd195;  #10 
a = 8'd152; b = 8'd196;  #10 
a = 8'd152; b = 8'd197;  #10 
a = 8'd152; b = 8'd198;  #10 
a = 8'd152; b = 8'd199;  #10 
a = 8'd152; b = 8'd200;  #10 
a = 8'd152; b = 8'd201;  #10 
a = 8'd152; b = 8'd202;  #10 
a = 8'd152; b = 8'd203;  #10 
a = 8'd152; b = 8'd204;  #10 
a = 8'd152; b = 8'd205;  #10 
a = 8'd152; b = 8'd206;  #10 
a = 8'd152; b = 8'd207;  #10 
a = 8'd152; b = 8'd208;  #10 
a = 8'd152; b = 8'd209;  #10 
a = 8'd152; b = 8'd210;  #10 
a = 8'd152; b = 8'd211;  #10 
a = 8'd152; b = 8'd212;  #10 
a = 8'd152; b = 8'd213;  #10 
a = 8'd152; b = 8'd214;  #10 
a = 8'd152; b = 8'd215;  #10 
a = 8'd152; b = 8'd216;  #10 
a = 8'd152; b = 8'd217;  #10 
a = 8'd152; b = 8'd218;  #10 
a = 8'd152; b = 8'd219;  #10 
a = 8'd152; b = 8'd220;  #10 
a = 8'd152; b = 8'd221;  #10 
a = 8'd152; b = 8'd222;  #10 
a = 8'd152; b = 8'd223;  #10 
a = 8'd152; b = 8'd224;  #10 
a = 8'd152; b = 8'd225;  #10 
a = 8'd152; b = 8'd226;  #10 
a = 8'd152; b = 8'd227;  #10 
a = 8'd152; b = 8'd228;  #10 
a = 8'd152; b = 8'd229;  #10 
a = 8'd152; b = 8'd230;  #10 
a = 8'd152; b = 8'd231;  #10 
a = 8'd152; b = 8'd232;  #10 
a = 8'd152; b = 8'd233;  #10 
a = 8'd152; b = 8'd234;  #10 
a = 8'd152; b = 8'd235;  #10 
a = 8'd152; b = 8'd236;  #10 
a = 8'd152; b = 8'd237;  #10 
a = 8'd152; b = 8'd238;  #10 
a = 8'd152; b = 8'd239;  #10 
a = 8'd152; b = 8'd240;  #10 
a = 8'd152; b = 8'd241;  #10 
a = 8'd152; b = 8'd242;  #10 
a = 8'd152; b = 8'd243;  #10 
a = 8'd152; b = 8'd244;  #10 
a = 8'd152; b = 8'd245;  #10 
a = 8'd152; b = 8'd246;  #10 
a = 8'd152; b = 8'd247;  #10 
a = 8'd152; b = 8'd248;  #10 
a = 8'd152; b = 8'd249;  #10 
a = 8'd152; b = 8'd250;  #10 
a = 8'd152; b = 8'd251;  #10 
a = 8'd152; b = 8'd252;  #10 
a = 8'd152; b = 8'd253;  #10 
a = 8'd152; b = 8'd254;  #10 
a = 8'd152; b = 8'd255;  #10 
a = 8'd153; b = 8'd0;  #10 
a = 8'd153; b = 8'd1;  #10 
a = 8'd153; b = 8'd2;  #10 
a = 8'd153; b = 8'd3;  #10 
a = 8'd153; b = 8'd4;  #10 
a = 8'd153; b = 8'd5;  #10 
a = 8'd153; b = 8'd6;  #10 
a = 8'd153; b = 8'd7;  #10 
a = 8'd153; b = 8'd8;  #10 
a = 8'd153; b = 8'd9;  #10 
a = 8'd153; b = 8'd10;  #10 
a = 8'd153; b = 8'd11;  #10 
a = 8'd153; b = 8'd12;  #10 
a = 8'd153; b = 8'd13;  #10 
a = 8'd153; b = 8'd14;  #10 
a = 8'd153; b = 8'd15;  #10 
a = 8'd153; b = 8'd16;  #10 
a = 8'd153; b = 8'd17;  #10 
a = 8'd153; b = 8'd18;  #10 
a = 8'd153; b = 8'd19;  #10 
a = 8'd153; b = 8'd20;  #10 
a = 8'd153; b = 8'd21;  #10 
a = 8'd153; b = 8'd22;  #10 
a = 8'd153; b = 8'd23;  #10 
a = 8'd153; b = 8'd24;  #10 
a = 8'd153; b = 8'd25;  #10 
a = 8'd153; b = 8'd26;  #10 
a = 8'd153; b = 8'd27;  #10 
a = 8'd153; b = 8'd28;  #10 
a = 8'd153; b = 8'd29;  #10 
a = 8'd153; b = 8'd30;  #10 
a = 8'd153; b = 8'd31;  #10 
a = 8'd153; b = 8'd32;  #10 
a = 8'd153; b = 8'd33;  #10 
a = 8'd153; b = 8'd34;  #10 
a = 8'd153; b = 8'd35;  #10 
a = 8'd153; b = 8'd36;  #10 
a = 8'd153; b = 8'd37;  #10 
a = 8'd153; b = 8'd38;  #10 
a = 8'd153; b = 8'd39;  #10 
a = 8'd153; b = 8'd40;  #10 
a = 8'd153; b = 8'd41;  #10 
a = 8'd153; b = 8'd42;  #10 
a = 8'd153; b = 8'd43;  #10 
a = 8'd153; b = 8'd44;  #10 
a = 8'd153; b = 8'd45;  #10 
a = 8'd153; b = 8'd46;  #10 
a = 8'd153; b = 8'd47;  #10 
a = 8'd153; b = 8'd48;  #10 
a = 8'd153; b = 8'd49;  #10 
a = 8'd153; b = 8'd50;  #10 
a = 8'd153; b = 8'd51;  #10 
a = 8'd153; b = 8'd52;  #10 
a = 8'd153; b = 8'd53;  #10 
a = 8'd153; b = 8'd54;  #10 
a = 8'd153; b = 8'd55;  #10 
a = 8'd153; b = 8'd56;  #10 
a = 8'd153; b = 8'd57;  #10 
a = 8'd153; b = 8'd58;  #10 
a = 8'd153; b = 8'd59;  #10 
a = 8'd153; b = 8'd60;  #10 
a = 8'd153; b = 8'd61;  #10 
a = 8'd153; b = 8'd62;  #10 
a = 8'd153; b = 8'd63;  #10 
a = 8'd153; b = 8'd64;  #10 
a = 8'd153; b = 8'd65;  #10 
a = 8'd153; b = 8'd66;  #10 
a = 8'd153; b = 8'd67;  #10 
a = 8'd153; b = 8'd68;  #10 
a = 8'd153; b = 8'd69;  #10 
a = 8'd153; b = 8'd70;  #10 
a = 8'd153; b = 8'd71;  #10 
a = 8'd153; b = 8'd72;  #10 
a = 8'd153; b = 8'd73;  #10 
a = 8'd153; b = 8'd74;  #10 
a = 8'd153; b = 8'd75;  #10 
a = 8'd153; b = 8'd76;  #10 
a = 8'd153; b = 8'd77;  #10 
a = 8'd153; b = 8'd78;  #10 
a = 8'd153; b = 8'd79;  #10 
a = 8'd153; b = 8'd80;  #10 
a = 8'd153; b = 8'd81;  #10 
a = 8'd153; b = 8'd82;  #10 
a = 8'd153; b = 8'd83;  #10 
a = 8'd153; b = 8'd84;  #10 
a = 8'd153; b = 8'd85;  #10 
a = 8'd153; b = 8'd86;  #10 
a = 8'd153; b = 8'd87;  #10 
a = 8'd153; b = 8'd88;  #10 
a = 8'd153; b = 8'd89;  #10 
a = 8'd153; b = 8'd90;  #10 
a = 8'd153; b = 8'd91;  #10 
a = 8'd153; b = 8'd92;  #10 
a = 8'd153; b = 8'd93;  #10 
a = 8'd153; b = 8'd94;  #10 
a = 8'd153; b = 8'd95;  #10 
a = 8'd153; b = 8'd96;  #10 
a = 8'd153; b = 8'd97;  #10 
a = 8'd153; b = 8'd98;  #10 
a = 8'd153; b = 8'd99;  #10 
a = 8'd153; b = 8'd100;  #10 
a = 8'd153; b = 8'd101;  #10 
a = 8'd153; b = 8'd102;  #10 
a = 8'd153; b = 8'd103;  #10 
a = 8'd153; b = 8'd104;  #10 
a = 8'd153; b = 8'd105;  #10 
a = 8'd153; b = 8'd106;  #10 
a = 8'd153; b = 8'd107;  #10 
a = 8'd153; b = 8'd108;  #10 
a = 8'd153; b = 8'd109;  #10 
a = 8'd153; b = 8'd110;  #10 
a = 8'd153; b = 8'd111;  #10 
a = 8'd153; b = 8'd112;  #10 
a = 8'd153; b = 8'd113;  #10 
a = 8'd153; b = 8'd114;  #10 
a = 8'd153; b = 8'd115;  #10 
a = 8'd153; b = 8'd116;  #10 
a = 8'd153; b = 8'd117;  #10 
a = 8'd153; b = 8'd118;  #10 
a = 8'd153; b = 8'd119;  #10 
a = 8'd153; b = 8'd120;  #10 
a = 8'd153; b = 8'd121;  #10 
a = 8'd153; b = 8'd122;  #10 
a = 8'd153; b = 8'd123;  #10 
a = 8'd153; b = 8'd124;  #10 
a = 8'd153; b = 8'd125;  #10 
a = 8'd153; b = 8'd126;  #10 
a = 8'd153; b = 8'd127;  #10 
a = 8'd153; b = 8'd128;  #10 
a = 8'd153; b = 8'd129;  #10 
a = 8'd153; b = 8'd130;  #10 
a = 8'd153; b = 8'd131;  #10 
a = 8'd153; b = 8'd132;  #10 
a = 8'd153; b = 8'd133;  #10 
a = 8'd153; b = 8'd134;  #10 
a = 8'd153; b = 8'd135;  #10 
a = 8'd153; b = 8'd136;  #10 
a = 8'd153; b = 8'd137;  #10 
a = 8'd153; b = 8'd138;  #10 
a = 8'd153; b = 8'd139;  #10 
a = 8'd153; b = 8'd140;  #10 
a = 8'd153; b = 8'd141;  #10 
a = 8'd153; b = 8'd142;  #10 
a = 8'd153; b = 8'd143;  #10 
a = 8'd153; b = 8'd144;  #10 
a = 8'd153; b = 8'd145;  #10 
a = 8'd153; b = 8'd146;  #10 
a = 8'd153; b = 8'd147;  #10 
a = 8'd153; b = 8'd148;  #10 
a = 8'd153; b = 8'd149;  #10 
a = 8'd153; b = 8'd150;  #10 
a = 8'd153; b = 8'd151;  #10 
a = 8'd153; b = 8'd152;  #10 
a = 8'd153; b = 8'd153;  #10 
a = 8'd153; b = 8'd154;  #10 
a = 8'd153; b = 8'd155;  #10 
a = 8'd153; b = 8'd156;  #10 
a = 8'd153; b = 8'd157;  #10 
a = 8'd153; b = 8'd158;  #10 
a = 8'd153; b = 8'd159;  #10 
a = 8'd153; b = 8'd160;  #10 
a = 8'd153; b = 8'd161;  #10 
a = 8'd153; b = 8'd162;  #10 
a = 8'd153; b = 8'd163;  #10 
a = 8'd153; b = 8'd164;  #10 
a = 8'd153; b = 8'd165;  #10 
a = 8'd153; b = 8'd166;  #10 
a = 8'd153; b = 8'd167;  #10 
a = 8'd153; b = 8'd168;  #10 
a = 8'd153; b = 8'd169;  #10 
a = 8'd153; b = 8'd170;  #10 
a = 8'd153; b = 8'd171;  #10 
a = 8'd153; b = 8'd172;  #10 
a = 8'd153; b = 8'd173;  #10 
a = 8'd153; b = 8'd174;  #10 
a = 8'd153; b = 8'd175;  #10 
a = 8'd153; b = 8'd176;  #10 
a = 8'd153; b = 8'd177;  #10 
a = 8'd153; b = 8'd178;  #10 
a = 8'd153; b = 8'd179;  #10 
a = 8'd153; b = 8'd180;  #10 
a = 8'd153; b = 8'd181;  #10 
a = 8'd153; b = 8'd182;  #10 
a = 8'd153; b = 8'd183;  #10 
a = 8'd153; b = 8'd184;  #10 
a = 8'd153; b = 8'd185;  #10 
a = 8'd153; b = 8'd186;  #10 
a = 8'd153; b = 8'd187;  #10 
a = 8'd153; b = 8'd188;  #10 
a = 8'd153; b = 8'd189;  #10 
a = 8'd153; b = 8'd190;  #10 
a = 8'd153; b = 8'd191;  #10 
a = 8'd153; b = 8'd192;  #10 
a = 8'd153; b = 8'd193;  #10 
a = 8'd153; b = 8'd194;  #10 
a = 8'd153; b = 8'd195;  #10 
a = 8'd153; b = 8'd196;  #10 
a = 8'd153; b = 8'd197;  #10 
a = 8'd153; b = 8'd198;  #10 
a = 8'd153; b = 8'd199;  #10 
a = 8'd153; b = 8'd200;  #10 
a = 8'd153; b = 8'd201;  #10 
a = 8'd153; b = 8'd202;  #10 
a = 8'd153; b = 8'd203;  #10 
a = 8'd153; b = 8'd204;  #10 
a = 8'd153; b = 8'd205;  #10 
a = 8'd153; b = 8'd206;  #10 
a = 8'd153; b = 8'd207;  #10 
a = 8'd153; b = 8'd208;  #10 
a = 8'd153; b = 8'd209;  #10 
a = 8'd153; b = 8'd210;  #10 
a = 8'd153; b = 8'd211;  #10 
a = 8'd153; b = 8'd212;  #10 
a = 8'd153; b = 8'd213;  #10 
a = 8'd153; b = 8'd214;  #10 
a = 8'd153; b = 8'd215;  #10 
a = 8'd153; b = 8'd216;  #10 
a = 8'd153; b = 8'd217;  #10 
a = 8'd153; b = 8'd218;  #10 
a = 8'd153; b = 8'd219;  #10 
a = 8'd153; b = 8'd220;  #10 
a = 8'd153; b = 8'd221;  #10 
a = 8'd153; b = 8'd222;  #10 
a = 8'd153; b = 8'd223;  #10 
a = 8'd153; b = 8'd224;  #10 
a = 8'd153; b = 8'd225;  #10 
a = 8'd153; b = 8'd226;  #10 
a = 8'd153; b = 8'd227;  #10 
a = 8'd153; b = 8'd228;  #10 
a = 8'd153; b = 8'd229;  #10 
a = 8'd153; b = 8'd230;  #10 
a = 8'd153; b = 8'd231;  #10 
a = 8'd153; b = 8'd232;  #10 
a = 8'd153; b = 8'd233;  #10 
a = 8'd153; b = 8'd234;  #10 
a = 8'd153; b = 8'd235;  #10 
a = 8'd153; b = 8'd236;  #10 
a = 8'd153; b = 8'd237;  #10 
a = 8'd153; b = 8'd238;  #10 
a = 8'd153; b = 8'd239;  #10 
a = 8'd153; b = 8'd240;  #10 
a = 8'd153; b = 8'd241;  #10 
a = 8'd153; b = 8'd242;  #10 
a = 8'd153; b = 8'd243;  #10 
a = 8'd153; b = 8'd244;  #10 
a = 8'd153; b = 8'd245;  #10 
a = 8'd153; b = 8'd246;  #10 
a = 8'd153; b = 8'd247;  #10 
a = 8'd153; b = 8'd248;  #10 
a = 8'd153; b = 8'd249;  #10 
a = 8'd153; b = 8'd250;  #10 
a = 8'd153; b = 8'd251;  #10 
a = 8'd153; b = 8'd252;  #10 
a = 8'd153; b = 8'd253;  #10 
a = 8'd153; b = 8'd254;  #10 
a = 8'd153; b = 8'd255;  #10 
a = 8'd154; b = 8'd0;  #10 
a = 8'd154; b = 8'd1;  #10 
a = 8'd154; b = 8'd2;  #10 
a = 8'd154; b = 8'd3;  #10 
a = 8'd154; b = 8'd4;  #10 
a = 8'd154; b = 8'd5;  #10 
a = 8'd154; b = 8'd6;  #10 
a = 8'd154; b = 8'd7;  #10 
a = 8'd154; b = 8'd8;  #10 
a = 8'd154; b = 8'd9;  #10 
a = 8'd154; b = 8'd10;  #10 
a = 8'd154; b = 8'd11;  #10 
a = 8'd154; b = 8'd12;  #10 
a = 8'd154; b = 8'd13;  #10 
a = 8'd154; b = 8'd14;  #10 
a = 8'd154; b = 8'd15;  #10 
a = 8'd154; b = 8'd16;  #10 
a = 8'd154; b = 8'd17;  #10 
a = 8'd154; b = 8'd18;  #10 
a = 8'd154; b = 8'd19;  #10 
a = 8'd154; b = 8'd20;  #10 
a = 8'd154; b = 8'd21;  #10 
a = 8'd154; b = 8'd22;  #10 
a = 8'd154; b = 8'd23;  #10 
a = 8'd154; b = 8'd24;  #10 
a = 8'd154; b = 8'd25;  #10 
a = 8'd154; b = 8'd26;  #10 
a = 8'd154; b = 8'd27;  #10 
a = 8'd154; b = 8'd28;  #10 
a = 8'd154; b = 8'd29;  #10 
a = 8'd154; b = 8'd30;  #10 
a = 8'd154; b = 8'd31;  #10 
a = 8'd154; b = 8'd32;  #10 
a = 8'd154; b = 8'd33;  #10 
a = 8'd154; b = 8'd34;  #10 
a = 8'd154; b = 8'd35;  #10 
a = 8'd154; b = 8'd36;  #10 
a = 8'd154; b = 8'd37;  #10 
a = 8'd154; b = 8'd38;  #10 
a = 8'd154; b = 8'd39;  #10 
a = 8'd154; b = 8'd40;  #10 
a = 8'd154; b = 8'd41;  #10 
a = 8'd154; b = 8'd42;  #10 
a = 8'd154; b = 8'd43;  #10 
a = 8'd154; b = 8'd44;  #10 
a = 8'd154; b = 8'd45;  #10 
a = 8'd154; b = 8'd46;  #10 
a = 8'd154; b = 8'd47;  #10 
a = 8'd154; b = 8'd48;  #10 
a = 8'd154; b = 8'd49;  #10 
a = 8'd154; b = 8'd50;  #10 
a = 8'd154; b = 8'd51;  #10 
a = 8'd154; b = 8'd52;  #10 
a = 8'd154; b = 8'd53;  #10 
a = 8'd154; b = 8'd54;  #10 
a = 8'd154; b = 8'd55;  #10 
a = 8'd154; b = 8'd56;  #10 
a = 8'd154; b = 8'd57;  #10 
a = 8'd154; b = 8'd58;  #10 
a = 8'd154; b = 8'd59;  #10 
a = 8'd154; b = 8'd60;  #10 
a = 8'd154; b = 8'd61;  #10 
a = 8'd154; b = 8'd62;  #10 
a = 8'd154; b = 8'd63;  #10 
a = 8'd154; b = 8'd64;  #10 
a = 8'd154; b = 8'd65;  #10 
a = 8'd154; b = 8'd66;  #10 
a = 8'd154; b = 8'd67;  #10 
a = 8'd154; b = 8'd68;  #10 
a = 8'd154; b = 8'd69;  #10 
a = 8'd154; b = 8'd70;  #10 
a = 8'd154; b = 8'd71;  #10 
a = 8'd154; b = 8'd72;  #10 
a = 8'd154; b = 8'd73;  #10 
a = 8'd154; b = 8'd74;  #10 
a = 8'd154; b = 8'd75;  #10 
a = 8'd154; b = 8'd76;  #10 
a = 8'd154; b = 8'd77;  #10 
a = 8'd154; b = 8'd78;  #10 
a = 8'd154; b = 8'd79;  #10 
a = 8'd154; b = 8'd80;  #10 
a = 8'd154; b = 8'd81;  #10 
a = 8'd154; b = 8'd82;  #10 
a = 8'd154; b = 8'd83;  #10 
a = 8'd154; b = 8'd84;  #10 
a = 8'd154; b = 8'd85;  #10 
a = 8'd154; b = 8'd86;  #10 
a = 8'd154; b = 8'd87;  #10 
a = 8'd154; b = 8'd88;  #10 
a = 8'd154; b = 8'd89;  #10 
a = 8'd154; b = 8'd90;  #10 
a = 8'd154; b = 8'd91;  #10 
a = 8'd154; b = 8'd92;  #10 
a = 8'd154; b = 8'd93;  #10 
a = 8'd154; b = 8'd94;  #10 
a = 8'd154; b = 8'd95;  #10 
a = 8'd154; b = 8'd96;  #10 
a = 8'd154; b = 8'd97;  #10 
a = 8'd154; b = 8'd98;  #10 
a = 8'd154; b = 8'd99;  #10 
a = 8'd154; b = 8'd100;  #10 
a = 8'd154; b = 8'd101;  #10 
a = 8'd154; b = 8'd102;  #10 
a = 8'd154; b = 8'd103;  #10 
a = 8'd154; b = 8'd104;  #10 
a = 8'd154; b = 8'd105;  #10 
a = 8'd154; b = 8'd106;  #10 
a = 8'd154; b = 8'd107;  #10 
a = 8'd154; b = 8'd108;  #10 
a = 8'd154; b = 8'd109;  #10 
a = 8'd154; b = 8'd110;  #10 
a = 8'd154; b = 8'd111;  #10 
a = 8'd154; b = 8'd112;  #10 
a = 8'd154; b = 8'd113;  #10 
a = 8'd154; b = 8'd114;  #10 
a = 8'd154; b = 8'd115;  #10 
a = 8'd154; b = 8'd116;  #10 
a = 8'd154; b = 8'd117;  #10 
a = 8'd154; b = 8'd118;  #10 
a = 8'd154; b = 8'd119;  #10 
a = 8'd154; b = 8'd120;  #10 
a = 8'd154; b = 8'd121;  #10 
a = 8'd154; b = 8'd122;  #10 
a = 8'd154; b = 8'd123;  #10 
a = 8'd154; b = 8'd124;  #10 
a = 8'd154; b = 8'd125;  #10 
a = 8'd154; b = 8'd126;  #10 
a = 8'd154; b = 8'd127;  #10 
a = 8'd154; b = 8'd128;  #10 
a = 8'd154; b = 8'd129;  #10 
a = 8'd154; b = 8'd130;  #10 
a = 8'd154; b = 8'd131;  #10 
a = 8'd154; b = 8'd132;  #10 
a = 8'd154; b = 8'd133;  #10 
a = 8'd154; b = 8'd134;  #10 
a = 8'd154; b = 8'd135;  #10 
a = 8'd154; b = 8'd136;  #10 
a = 8'd154; b = 8'd137;  #10 
a = 8'd154; b = 8'd138;  #10 
a = 8'd154; b = 8'd139;  #10 
a = 8'd154; b = 8'd140;  #10 
a = 8'd154; b = 8'd141;  #10 
a = 8'd154; b = 8'd142;  #10 
a = 8'd154; b = 8'd143;  #10 
a = 8'd154; b = 8'd144;  #10 
a = 8'd154; b = 8'd145;  #10 
a = 8'd154; b = 8'd146;  #10 
a = 8'd154; b = 8'd147;  #10 
a = 8'd154; b = 8'd148;  #10 
a = 8'd154; b = 8'd149;  #10 
a = 8'd154; b = 8'd150;  #10 
a = 8'd154; b = 8'd151;  #10 
a = 8'd154; b = 8'd152;  #10 
a = 8'd154; b = 8'd153;  #10 
a = 8'd154; b = 8'd154;  #10 
a = 8'd154; b = 8'd155;  #10 
a = 8'd154; b = 8'd156;  #10 
a = 8'd154; b = 8'd157;  #10 
a = 8'd154; b = 8'd158;  #10 
a = 8'd154; b = 8'd159;  #10 
a = 8'd154; b = 8'd160;  #10 
a = 8'd154; b = 8'd161;  #10 
a = 8'd154; b = 8'd162;  #10 
a = 8'd154; b = 8'd163;  #10 
a = 8'd154; b = 8'd164;  #10 
a = 8'd154; b = 8'd165;  #10 
a = 8'd154; b = 8'd166;  #10 
a = 8'd154; b = 8'd167;  #10 
a = 8'd154; b = 8'd168;  #10 
a = 8'd154; b = 8'd169;  #10 
a = 8'd154; b = 8'd170;  #10 
a = 8'd154; b = 8'd171;  #10 
a = 8'd154; b = 8'd172;  #10 
a = 8'd154; b = 8'd173;  #10 
a = 8'd154; b = 8'd174;  #10 
a = 8'd154; b = 8'd175;  #10 
a = 8'd154; b = 8'd176;  #10 
a = 8'd154; b = 8'd177;  #10 
a = 8'd154; b = 8'd178;  #10 
a = 8'd154; b = 8'd179;  #10 
a = 8'd154; b = 8'd180;  #10 
a = 8'd154; b = 8'd181;  #10 
a = 8'd154; b = 8'd182;  #10 
a = 8'd154; b = 8'd183;  #10 
a = 8'd154; b = 8'd184;  #10 
a = 8'd154; b = 8'd185;  #10 
a = 8'd154; b = 8'd186;  #10 
a = 8'd154; b = 8'd187;  #10 
a = 8'd154; b = 8'd188;  #10 
a = 8'd154; b = 8'd189;  #10 
a = 8'd154; b = 8'd190;  #10 
a = 8'd154; b = 8'd191;  #10 
a = 8'd154; b = 8'd192;  #10 
a = 8'd154; b = 8'd193;  #10 
a = 8'd154; b = 8'd194;  #10 
a = 8'd154; b = 8'd195;  #10 
a = 8'd154; b = 8'd196;  #10 
a = 8'd154; b = 8'd197;  #10 
a = 8'd154; b = 8'd198;  #10 
a = 8'd154; b = 8'd199;  #10 
a = 8'd154; b = 8'd200;  #10 
a = 8'd154; b = 8'd201;  #10 
a = 8'd154; b = 8'd202;  #10 
a = 8'd154; b = 8'd203;  #10 
a = 8'd154; b = 8'd204;  #10 
a = 8'd154; b = 8'd205;  #10 
a = 8'd154; b = 8'd206;  #10 
a = 8'd154; b = 8'd207;  #10 
a = 8'd154; b = 8'd208;  #10 
a = 8'd154; b = 8'd209;  #10 
a = 8'd154; b = 8'd210;  #10 
a = 8'd154; b = 8'd211;  #10 
a = 8'd154; b = 8'd212;  #10 
a = 8'd154; b = 8'd213;  #10 
a = 8'd154; b = 8'd214;  #10 
a = 8'd154; b = 8'd215;  #10 
a = 8'd154; b = 8'd216;  #10 
a = 8'd154; b = 8'd217;  #10 
a = 8'd154; b = 8'd218;  #10 
a = 8'd154; b = 8'd219;  #10 
a = 8'd154; b = 8'd220;  #10 
a = 8'd154; b = 8'd221;  #10 
a = 8'd154; b = 8'd222;  #10 
a = 8'd154; b = 8'd223;  #10 
a = 8'd154; b = 8'd224;  #10 
a = 8'd154; b = 8'd225;  #10 
a = 8'd154; b = 8'd226;  #10 
a = 8'd154; b = 8'd227;  #10 
a = 8'd154; b = 8'd228;  #10 
a = 8'd154; b = 8'd229;  #10 
a = 8'd154; b = 8'd230;  #10 
a = 8'd154; b = 8'd231;  #10 
a = 8'd154; b = 8'd232;  #10 
a = 8'd154; b = 8'd233;  #10 
a = 8'd154; b = 8'd234;  #10 
a = 8'd154; b = 8'd235;  #10 
a = 8'd154; b = 8'd236;  #10 
a = 8'd154; b = 8'd237;  #10 
a = 8'd154; b = 8'd238;  #10 
a = 8'd154; b = 8'd239;  #10 
a = 8'd154; b = 8'd240;  #10 
a = 8'd154; b = 8'd241;  #10 
a = 8'd154; b = 8'd242;  #10 
a = 8'd154; b = 8'd243;  #10 
a = 8'd154; b = 8'd244;  #10 
a = 8'd154; b = 8'd245;  #10 
a = 8'd154; b = 8'd246;  #10 
a = 8'd154; b = 8'd247;  #10 
a = 8'd154; b = 8'd248;  #10 
a = 8'd154; b = 8'd249;  #10 
a = 8'd154; b = 8'd250;  #10 
a = 8'd154; b = 8'd251;  #10 
a = 8'd154; b = 8'd252;  #10 
a = 8'd154; b = 8'd253;  #10 
a = 8'd154; b = 8'd254;  #10 
a = 8'd154; b = 8'd255;  #10 
a = 8'd155; b = 8'd0;  #10 
a = 8'd155; b = 8'd1;  #10 
a = 8'd155; b = 8'd2;  #10 
a = 8'd155; b = 8'd3;  #10 
a = 8'd155; b = 8'd4;  #10 
a = 8'd155; b = 8'd5;  #10 
a = 8'd155; b = 8'd6;  #10 
a = 8'd155; b = 8'd7;  #10 
a = 8'd155; b = 8'd8;  #10 
a = 8'd155; b = 8'd9;  #10 
a = 8'd155; b = 8'd10;  #10 
a = 8'd155; b = 8'd11;  #10 
a = 8'd155; b = 8'd12;  #10 
a = 8'd155; b = 8'd13;  #10 
a = 8'd155; b = 8'd14;  #10 
a = 8'd155; b = 8'd15;  #10 
a = 8'd155; b = 8'd16;  #10 
a = 8'd155; b = 8'd17;  #10 
a = 8'd155; b = 8'd18;  #10 
a = 8'd155; b = 8'd19;  #10 
a = 8'd155; b = 8'd20;  #10 
a = 8'd155; b = 8'd21;  #10 
a = 8'd155; b = 8'd22;  #10 
a = 8'd155; b = 8'd23;  #10 
a = 8'd155; b = 8'd24;  #10 
a = 8'd155; b = 8'd25;  #10 
a = 8'd155; b = 8'd26;  #10 
a = 8'd155; b = 8'd27;  #10 
a = 8'd155; b = 8'd28;  #10 
a = 8'd155; b = 8'd29;  #10 
a = 8'd155; b = 8'd30;  #10 
a = 8'd155; b = 8'd31;  #10 
a = 8'd155; b = 8'd32;  #10 
a = 8'd155; b = 8'd33;  #10 
a = 8'd155; b = 8'd34;  #10 
a = 8'd155; b = 8'd35;  #10 
a = 8'd155; b = 8'd36;  #10 
a = 8'd155; b = 8'd37;  #10 
a = 8'd155; b = 8'd38;  #10 
a = 8'd155; b = 8'd39;  #10 
a = 8'd155; b = 8'd40;  #10 
a = 8'd155; b = 8'd41;  #10 
a = 8'd155; b = 8'd42;  #10 
a = 8'd155; b = 8'd43;  #10 
a = 8'd155; b = 8'd44;  #10 
a = 8'd155; b = 8'd45;  #10 
a = 8'd155; b = 8'd46;  #10 
a = 8'd155; b = 8'd47;  #10 
a = 8'd155; b = 8'd48;  #10 
a = 8'd155; b = 8'd49;  #10 
a = 8'd155; b = 8'd50;  #10 
a = 8'd155; b = 8'd51;  #10 
a = 8'd155; b = 8'd52;  #10 
a = 8'd155; b = 8'd53;  #10 
a = 8'd155; b = 8'd54;  #10 
a = 8'd155; b = 8'd55;  #10 
a = 8'd155; b = 8'd56;  #10 
a = 8'd155; b = 8'd57;  #10 
a = 8'd155; b = 8'd58;  #10 
a = 8'd155; b = 8'd59;  #10 
a = 8'd155; b = 8'd60;  #10 
a = 8'd155; b = 8'd61;  #10 
a = 8'd155; b = 8'd62;  #10 
a = 8'd155; b = 8'd63;  #10 
a = 8'd155; b = 8'd64;  #10 
a = 8'd155; b = 8'd65;  #10 
a = 8'd155; b = 8'd66;  #10 
a = 8'd155; b = 8'd67;  #10 
a = 8'd155; b = 8'd68;  #10 
a = 8'd155; b = 8'd69;  #10 
a = 8'd155; b = 8'd70;  #10 
a = 8'd155; b = 8'd71;  #10 
a = 8'd155; b = 8'd72;  #10 
a = 8'd155; b = 8'd73;  #10 
a = 8'd155; b = 8'd74;  #10 
a = 8'd155; b = 8'd75;  #10 
a = 8'd155; b = 8'd76;  #10 
a = 8'd155; b = 8'd77;  #10 
a = 8'd155; b = 8'd78;  #10 
a = 8'd155; b = 8'd79;  #10 
a = 8'd155; b = 8'd80;  #10 
a = 8'd155; b = 8'd81;  #10 
a = 8'd155; b = 8'd82;  #10 
a = 8'd155; b = 8'd83;  #10 
a = 8'd155; b = 8'd84;  #10 
a = 8'd155; b = 8'd85;  #10 
a = 8'd155; b = 8'd86;  #10 
a = 8'd155; b = 8'd87;  #10 
a = 8'd155; b = 8'd88;  #10 
a = 8'd155; b = 8'd89;  #10 
a = 8'd155; b = 8'd90;  #10 
a = 8'd155; b = 8'd91;  #10 
a = 8'd155; b = 8'd92;  #10 
a = 8'd155; b = 8'd93;  #10 
a = 8'd155; b = 8'd94;  #10 
a = 8'd155; b = 8'd95;  #10 
a = 8'd155; b = 8'd96;  #10 
a = 8'd155; b = 8'd97;  #10 
a = 8'd155; b = 8'd98;  #10 
a = 8'd155; b = 8'd99;  #10 
a = 8'd155; b = 8'd100;  #10 
a = 8'd155; b = 8'd101;  #10 
a = 8'd155; b = 8'd102;  #10 
a = 8'd155; b = 8'd103;  #10 
a = 8'd155; b = 8'd104;  #10 
a = 8'd155; b = 8'd105;  #10 
a = 8'd155; b = 8'd106;  #10 
a = 8'd155; b = 8'd107;  #10 
a = 8'd155; b = 8'd108;  #10 
a = 8'd155; b = 8'd109;  #10 
a = 8'd155; b = 8'd110;  #10 
a = 8'd155; b = 8'd111;  #10 
a = 8'd155; b = 8'd112;  #10 
a = 8'd155; b = 8'd113;  #10 
a = 8'd155; b = 8'd114;  #10 
a = 8'd155; b = 8'd115;  #10 
a = 8'd155; b = 8'd116;  #10 
a = 8'd155; b = 8'd117;  #10 
a = 8'd155; b = 8'd118;  #10 
a = 8'd155; b = 8'd119;  #10 
a = 8'd155; b = 8'd120;  #10 
a = 8'd155; b = 8'd121;  #10 
a = 8'd155; b = 8'd122;  #10 
a = 8'd155; b = 8'd123;  #10 
a = 8'd155; b = 8'd124;  #10 
a = 8'd155; b = 8'd125;  #10 
a = 8'd155; b = 8'd126;  #10 
a = 8'd155; b = 8'd127;  #10 
a = 8'd155; b = 8'd128;  #10 
a = 8'd155; b = 8'd129;  #10 
a = 8'd155; b = 8'd130;  #10 
a = 8'd155; b = 8'd131;  #10 
a = 8'd155; b = 8'd132;  #10 
a = 8'd155; b = 8'd133;  #10 
a = 8'd155; b = 8'd134;  #10 
a = 8'd155; b = 8'd135;  #10 
a = 8'd155; b = 8'd136;  #10 
a = 8'd155; b = 8'd137;  #10 
a = 8'd155; b = 8'd138;  #10 
a = 8'd155; b = 8'd139;  #10 
a = 8'd155; b = 8'd140;  #10 
a = 8'd155; b = 8'd141;  #10 
a = 8'd155; b = 8'd142;  #10 
a = 8'd155; b = 8'd143;  #10 
a = 8'd155; b = 8'd144;  #10 
a = 8'd155; b = 8'd145;  #10 
a = 8'd155; b = 8'd146;  #10 
a = 8'd155; b = 8'd147;  #10 
a = 8'd155; b = 8'd148;  #10 
a = 8'd155; b = 8'd149;  #10 
a = 8'd155; b = 8'd150;  #10 
a = 8'd155; b = 8'd151;  #10 
a = 8'd155; b = 8'd152;  #10 
a = 8'd155; b = 8'd153;  #10 
a = 8'd155; b = 8'd154;  #10 
a = 8'd155; b = 8'd155;  #10 
a = 8'd155; b = 8'd156;  #10 
a = 8'd155; b = 8'd157;  #10 
a = 8'd155; b = 8'd158;  #10 
a = 8'd155; b = 8'd159;  #10 
a = 8'd155; b = 8'd160;  #10 
a = 8'd155; b = 8'd161;  #10 
a = 8'd155; b = 8'd162;  #10 
a = 8'd155; b = 8'd163;  #10 
a = 8'd155; b = 8'd164;  #10 
a = 8'd155; b = 8'd165;  #10 
a = 8'd155; b = 8'd166;  #10 
a = 8'd155; b = 8'd167;  #10 
a = 8'd155; b = 8'd168;  #10 
a = 8'd155; b = 8'd169;  #10 
a = 8'd155; b = 8'd170;  #10 
a = 8'd155; b = 8'd171;  #10 
a = 8'd155; b = 8'd172;  #10 
a = 8'd155; b = 8'd173;  #10 
a = 8'd155; b = 8'd174;  #10 
a = 8'd155; b = 8'd175;  #10 
a = 8'd155; b = 8'd176;  #10 
a = 8'd155; b = 8'd177;  #10 
a = 8'd155; b = 8'd178;  #10 
a = 8'd155; b = 8'd179;  #10 
a = 8'd155; b = 8'd180;  #10 
a = 8'd155; b = 8'd181;  #10 
a = 8'd155; b = 8'd182;  #10 
a = 8'd155; b = 8'd183;  #10 
a = 8'd155; b = 8'd184;  #10 
a = 8'd155; b = 8'd185;  #10 
a = 8'd155; b = 8'd186;  #10 
a = 8'd155; b = 8'd187;  #10 
a = 8'd155; b = 8'd188;  #10 
a = 8'd155; b = 8'd189;  #10 
a = 8'd155; b = 8'd190;  #10 
a = 8'd155; b = 8'd191;  #10 
a = 8'd155; b = 8'd192;  #10 
a = 8'd155; b = 8'd193;  #10 
a = 8'd155; b = 8'd194;  #10 
a = 8'd155; b = 8'd195;  #10 
a = 8'd155; b = 8'd196;  #10 
a = 8'd155; b = 8'd197;  #10 
a = 8'd155; b = 8'd198;  #10 
a = 8'd155; b = 8'd199;  #10 
a = 8'd155; b = 8'd200;  #10 
a = 8'd155; b = 8'd201;  #10 
a = 8'd155; b = 8'd202;  #10 
a = 8'd155; b = 8'd203;  #10 
a = 8'd155; b = 8'd204;  #10 
a = 8'd155; b = 8'd205;  #10 
a = 8'd155; b = 8'd206;  #10 
a = 8'd155; b = 8'd207;  #10 
a = 8'd155; b = 8'd208;  #10 
a = 8'd155; b = 8'd209;  #10 
a = 8'd155; b = 8'd210;  #10 
a = 8'd155; b = 8'd211;  #10 
a = 8'd155; b = 8'd212;  #10 
a = 8'd155; b = 8'd213;  #10 
a = 8'd155; b = 8'd214;  #10 
a = 8'd155; b = 8'd215;  #10 
a = 8'd155; b = 8'd216;  #10 
a = 8'd155; b = 8'd217;  #10 
a = 8'd155; b = 8'd218;  #10 
a = 8'd155; b = 8'd219;  #10 
a = 8'd155; b = 8'd220;  #10 
a = 8'd155; b = 8'd221;  #10 
a = 8'd155; b = 8'd222;  #10 
a = 8'd155; b = 8'd223;  #10 
a = 8'd155; b = 8'd224;  #10 
a = 8'd155; b = 8'd225;  #10 
a = 8'd155; b = 8'd226;  #10 
a = 8'd155; b = 8'd227;  #10 
a = 8'd155; b = 8'd228;  #10 
a = 8'd155; b = 8'd229;  #10 
a = 8'd155; b = 8'd230;  #10 
a = 8'd155; b = 8'd231;  #10 
a = 8'd155; b = 8'd232;  #10 
a = 8'd155; b = 8'd233;  #10 
a = 8'd155; b = 8'd234;  #10 
a = 8'd155; b = 8'd235;  #10 
a = 8'd155; b = 8'd236;  #10 
a = 8'd155; b = 8'd237;  #10 
a = 8'd155; b = 8'd238;  #10 
a = 8'd155; b = 8'd239;  #10 
a = 8'd155; b = 8'd240;  #10 
a = 8'd155; b = 8'd241;  #10 
a = 8'd155; b = 8'd242;  #10 
a = 8'd155; b = 8'd243;  #10 
a = 8'd155; b = 8'd244;  #10 
a = 8'd155; b = 8'd245;  #10 
a = 8'd155; b = 8'd246;  #10 
a = 8'd155; b = 8'd247;  #10 
a = 8'd155; b = 8'd248;  #10 
a = 8'd155; b = 8'd249;  #10 
a = 8'd155; b = 8'd250;  #10 
a = 8'd155; b = 8'd251;  #10 
a = 8'd155; b = 8'd252;  #10 
a = 8'd155; b = 8'd253;  #10 
a = 8'd155; b = 8'd254;  #10 
a = 8'd155; b = 8'd255;  #10 
a = 8'd156; b = 8'd0;  #10 
a = 8'd156; b = 8'd1;  #10 
a = 8'd156; b = 8'd2;  #10 
a = 8'd156; b = 8'd3;  #10 
a = 8'd156; b = 8'd4;  #10 
a = 8'd156; b = 8'd5;  #10 
a = 8'd156; b = 8'd6;  #10 
a = 8'd156; b = 8'd7;  #10 
a = 8'd156; b = 8'd8;  #10 
a = 8'd156; b = 8'd9;  #10 
a = 8'd156; b = 8'd10;  #10 
a = 8'd156; b = 8'd11;  #10 
a = 8'd156; b = 8'd12;  #10 
a = 8'd156; b = 8'd13;  #10 
a = 8'd156; b = 8'd14;  #10 
a = 8'd156; b = 8'd15;  #10 
a = 8'd156; b = 8'd16;  #10 
a = 8'd156; b = 8'd17;  #10 
a = 8'd156; b = 8'd18;  #10 
a = 8'd156; b = 8'd19;  #10 
a = 8'd156; b = 8'd20;  #10 
a = 8'd156; b = 8'd21;  #10 
a = 8'd156; b = 8'd22;  #10 
a = 8'd156; b = 8'd23;  #10 
a = 8'd156; b = 8'd24;  #10 
a = 8'd156; b = 8'd25;  #10 
a = 8'd156; b = 8'd26;  #10 
a = 8'd156; b = 8'd27;  #10 
a = 8'd156; b = 8'd28;  #10 
a = 8'd156; b = 8'd29;  #10 
a = 8'd156; b = 8'd30;  #10 
a = 8'd156; b = 8'd31;  #10 
a = 8'd156; b = 8'd32;  #10 
a = 8'd156; b = 8'd33;  #10 
a = 8'd156; b = 8'd34;  #10 
a = 8'd156; b = 8'd35;  #10 
a = 8'd156; b = 8'd36;  #10 
a = 8'd156; b = 8'd37;  #10 
a = 8'd156; b = 8'd38;  #10 
a = 8'd156; b = 8'd39;  #10 
a = 8'd156; b = 8'd40;  #10 
a = 8'd156; b = 8'd41;  #10 
a = 8'd156; b = 8'd42;  #10 
a = 8'd156; b = 8'd43;  #10 
a = 8'd156; b = 8'd44;  #10 
a = 8'd156; b = 8'd45;  #10 
a = 8'd156; b = 8'd46;  #10 
a = 8'd156; b = 8'd47;  #10 
a = 8'd156; b = 8'd48;  #10 
a = 8'd156; b = 8'd49;  #10 
a = 8'd156; b = 8'd50;  #10 
a = 8'd156; b = 8'd51;  #10 
a = 8'd156; b = 8'd52;  #10 
a = 8'd156; b = 8'd53;  #10 
a = 8'd156; b = 8'd54;  #10 
a = 8'd156; b = 8'd55;  #10 
a = 8'd156; b = 8'd56;  #10 
a = 8'd156; b = 8'd57;  #10 
a = 8'd156; b = 8'd58;  #10 
a = 8'd156; b = 8'd59;  #10 
a = 8'd156; b = 8'd60;  #10 
a = 8'd156; b = 8'd61;  #10 
a = 8'd156; b = 8'd62;  #10 
a = 8'd156; b = 8'd63;  #10 
a = 8'd156; b = 8'd64;  #10 
a = 8'd156; b = 8'd65;  #10 
a = 8'd156; b = 8'd66;  #10 
a = 8'd156; b = 8'd67;  #10 
a = 8'd156; b = 8'd68;  #10 
a = 8'd156; b = 8'd69;  #10 
a = 8'd156; b = 8'd70;  #10 
a = 8'd156; b = 8'd71;  #10 
a = 8'd156; b = 8'd72;  #10 
a = 8'd156; b = 8'd73;  #10 
a = 8'd156; b = 8'd74;  #10 
a = 8'd156; b = 8'd75;  #10 
a = 8'd156; b = 8'd76;  #10 
a = 8'd156; b = 8'd77;  #10 
a = 8'd156; b = 8'd78;  #10 
a = 8'd156; b = 8'd79;  #10 
a = 8'd156; b = 8'd80;  #10 
a = 8'd156; b = 8'd81;  #10 
a = 8'd156; b = 8'd82;  #10 
a = 8'd156; b = 8'd83;  #10 
a = 8'd156; b = 8'd84;  #10 
a = 8'd156; b = 8'd85;  #10 
a = 8'd156; b = 8'd86;  #10 
a = 8'd156; b = 8'd87;  #10 
a = 8'd156; b = 8'd88;  #10 
a = 8'd156; b = 8'd89;  #10 
a = 8'd156; b = 8'd90;  #10 
a = 8'd156; b = 8'd91;  #10 
a = 8'd156; b = 8'd92;  #10 
a = 8'd156; b = 8'd93;  #10 
a = 8'd156; b = 8'd94;  #10 
a = 8'd156; b = 8'd95;  #10 
a = 8'd156; b = 8'd96;  #10 
a = 8'd156; b = 8'd97;  #10 
a = 8'd156; b = 8'd98;  #10 
a = 8'd156; b = 8'd99;  #10 
a = 8'd156; b = 8'd100;  #10 
a = 8'd156; b = 8'd101;  #10 
a = 8'd156; b = 8'd102;  #10 
a = 8'd156; b = 8'd103;  #10 
a = 8'd156; b = 8'd104;  #10 
a = 8'd156; b = 8'd105;  #10 
a = 8'd156; b = 8'd106;  #10 
a = 8'd156; b = 8'd107;  #10 
a = 8'd156; b = 8'd108;  #10 
a = 8'd156; b = 8'd109;  #10 
a = 8'd156; b = 8'd110;  #10 
a = 8'd156; b = 8'd111;  #10 
a = 8'd156; b = 8'd112;  #10 
a = 8'd156; b = 8'd113;  #10 
a = 8'd156; b = 8'd114;  #10 
a = 8'd156; b = 8'd115;  #10 
a = 8'd156; b = 8'd116;  #10 
a = 8'd156; b = 8'd117;  #10 
a = 8'd156; b = 8'd118;  #10 
a = 8'd156; b = 8'd119;  #10 
a = 8'd156; b = 8'd120;  #10 
a = 8'd156; b = 8'd121;  #10 
a = 8'd156; b = 8'd122;  #10 
a = 8'd156; b = 8'd123;  #10 
a = 8'd156; b = 8'd124;  #10 
a = 8'd156; b = 8'd125;  #10 
a = 8'd156; b = 8'd126;  #10 
a = 8'd156; b = 8'd127;  #10 
a = 8'd156; b = 8'd128;  #10 
a = 8'd156; b = 8'd129;  #10 
a = 8'd156; b = 8'd130;  #10 
a = 8'd156; b = 8'd131;  #10 
a = 8'd156; b = 8'd132;  #10 
a = 8'd156; b = 8'd133;  #10 
a = 8'd156; b = 8'd134;  #10 
a = 8'd156; b = 8'd135;  #10 
a = 8'd156; b = 8'd136;  #10 
a = 8'd156; b = 8'd137;  #10 
a = 8'd156; b = 8'd138;  #10 
a = 8'd156; b = 8'd139;  #10 
a = 8'd156; b = 8'd140;  #10 
a = 8'd156; b = 8'd141;  #10 
a = 8'd156; b = 8'd142;  #10 
a = 8'd156; b = 8'd143;  #10 
a = 8'd156; b = 8'd144;  #10 
a = 8'd156; b = 8'd145;  #10 
a = 8'd156; b = 8'd146;  #10 
a = 8'd156; b = 8'd147;  #10 
a = 8'd156; b = 8'd148;  #10 
a = 8'd156; b = 8'd149;  #10 
a = 8'd156; b = 8'd150;  #10 
a = 8'd156; b = 8'd151;  #10 
a = 8'd156; b = 8'd152;  #10 
a = 8'd156; b = 8'd153;  #10 
a = 8'd156; b = 8'd154;  #10 
a = 8'd156; b = 8'd155;  #10 
a = 8'd156; b = 8'd156;  #10 
a = 8'd156; b = 8'd157;  #10 
a = 8'd156; b = 8'd158;  #10 
a = 8'd156; b = 8'd159;  #10 
a = 8'd156; b = 8'd160;  #10 
a = 8'd156; b = 8'd161;  #10 
a = 8'd156; b = 8'd162;  #10 
a = 8'd156; b = 8'd163;  #10 
a = 8'd156; b = 8'd164;  #10 
a = 8'd156; b = 8'd165;  #10 
a = 8'd156; b = 8'd166;  #10 
a = 8'd156; b = 8'd167;  #10 
a = 8'd156; b = 8'd168;  #10 
a = 8'd156; b = 8'd169;  #10 
a = 8'd156; b = 8'd170;  #10 
a = 8'd156; b = 8'd171;  #10 
a = 8'd156; b = 8'd172;  #10 
a = 8'd156; b = 8'd173;  #10 
a = 8'd156; b = 8'd174;  #10 
a = 8'd156; b = 8'd175;  #10 
a = 8'd156; b = 8'd176;  #10 
a = 8'd156; b = 8'd177;  #10 
a = 8'd156; b = 8'd178;  #10 
a = 8'd156; b = 8'd179;  #10 
a = 8'd156; b = 8'd180;  #10 
a = 8'd156; b = 8'd181;  #10 
a = 8'd156; b = 8'd182;  #10 
a = 8'd156; b = 8'd183;  #10 
a = 8'd156; b = 8'd184;  #10 
a = 8'd156; b = 8'd185;  #10 
a = 8'd156; b = 8'd186;  #10 
a = 8'd156; b = 8'd187;  #10 
a = 8'd156; b = 8'd188;  #10 
a = 8'd156; b = 8'd189;  #10 
a = 8'd156; b = 8'd190;  #10 
a = 8'd156; b = 8'd191;  #10 
a = 8'd156; b = 8'd192;  #10 
a = 8'd156; b = 8'd193;  #10 
a = 8'd156; b = 8'd194;  #10 
a = 8'd156; b = 8'd195;  #10 
a = 8'd156; b = 8'd196;  #10 
a = 8'd156; b = 8'd197;  #10 
a = 8'd156; b = 8'd198;  #10 
a = 8'd156; b = 8'd199;  #10 
a = 8'd156; b = 8'd200;  #10 
a = 8'd156; b = 8'd201;  #10 
a = 8'd156; b = 8'd202;  #10 
a = 8'd156; b = 8'd203;  #10 
a = 8'd156; b = 8'd204;  #10 
a = 8'd156; b = 8'd205;  #10 
a = 8'd156; b = 8'd206;  #10 
a = 8'd156; b = 8'd207;  #10 
a = 8'd156; b = 8'd208;  #10 
a = 8'd156; b = 8'd209;  #10 
a = 8'd156; b = 8'd210;  #10 
a = 8'd156; b = 8'd211;  #10 
a = 8'd156; b = 8'd212;  #10 
a = 8'd156; b = 8'd213;  #10 
a = 8'd156; b = 8'd214;  #10 
a = 8'd156; b = 8'd215;  #10 
a = 8'd156; b = 8'd216;  #10 
a = 8'd156; b = 8'd217;  #10 
a = 8'd156; b = 8'd218;  #10 
a = 8'd156; b = 8'd219;  #10 
a = 8'd156; b = 8'd220;  #10 
a = 8'd156; b = 8'd221;  #10 
a = 8'd156; b = 8'd222;  #10 
a = 8'd156; b = 8'd223;  #10 
a = 8'd156; b = 8'd224;  #10 
a = 8'd156; b = 8'd225;  #10 
a = 8'd156; b = 8'd226;  #10 
a = 8'd156; b = 8'd227;  #10 
a = 8'd156; b = 8'd228;  #10 
a = 8'd156; b = 8'd229;  #10 
a = 8'd156; b = 8'd230;  #10 
a = 8'd156; b = 8'd231;  #10 
a = 8'd156; b = 8'd232;  #10 
a = 8'd156; b = 8'd233;  #10 
a = 8'd156; b = 8'd234;  #10 
a = 8'd156; b = 8'd235;  #10 
a = 8'd156; b = 8'd236;  #10 
a = 8'd156; b = 8'd237;  #10 
a = 8'd156; b = 8'd238;  #10 
a = 8'd156; b = 8'd239;  #10 
a = 8'd156; b = 8'd240;  #10 
a = 8'd156; b = 8'd241;  #10 
a = 8'd156; b = 8'd242;  #10 
a = 8'd156; b = 8'd243;  #10 
a = 8'd156; b = 8'd244;  #10 
a = 8'd156; b = 8'd245;  #10 
a = 8'd156; b = 8'd246;  #10 
a = 8'd156; b = 8'd247;  #10 
a = 8'd156; b = 8'd248;  #10 
a = 8'd156; b = 8'd249;  #10 
a = 8'd156; b = 8'd250;  #10 
a = 8'd156; b = 8'd251;  #10 
a = 8'd156; b = 8'd252;  #10 
a = 8'd156; b = 8'd253;  #10 
a = 8'd156; b = 8'd254;  #10 
a = 8'd156; b = 8'd255;  #10 
a = 8'd157; b = 8'd0;  #10 
a = 8'd157; b = 8'd1;  #10 
a = 8'd157; b = 8'd2;  #10 
a = 8'd157; b = 8'd3;  #10 
a = 8'd157; b = 8'd4;  #10 
a = 8'd157; b = 8'd5;  #10 
a = 8'd157; b = 8'd6;  #10 
a = 8'd157; b = 8'd7;  #10 
a = 8'd157; b = 8'd8;  #10 
a = 8'd157; b = 8'd9;  #10 
a = 8'd157; b = 8'd10;  #10 
a = 8'd157; b = 8'd11;  #10 
a = 8'd157; b = 8'd12;  #10 
a = 8'd157; b = 8'd13;  #10 
a = 8'd157; b = 8'd14;  #10 
a = 8'd157; b = 8'd15;  #10 
a = 8'd157; b = 8'd16;  #10 
a = 8'd157; b = 8'd17;  #10 
a = 8'd157; b = 8'd18;  #10 
a = 8'd157; b = 8'd19;  #10 
a = 8'd157; b = 8'd20;  #10 
a = 8'd157; b = 8'd21;  #10 
a = 8'd157; b = 8'd22;  #10 
a = 8'd157; b = 8'd23;  #10 
a = 8'd157; b = 8'd24;  #10 
a = 8'd157; b = 8'd25;  #10 
a = 8'd157; b = 8'd26;  #10 
a = 8'd157; b = 8'd27;  #10 
a = 8'd157; b = 8'd28;  #10 
a = 8'd157; b = 8'd29;  #10 
a = 8'd157; b = 8'd30;  #10 
a = 8'd157; b = 8'd31;  #10 
a = 8'd157; b = 8'd32;  #10 
a = 8'd157; b = 8'd33;  #10 
a = 8'd157; b = 8'd34;  #10 
a = 8'd157; b = 8'd35;  #10 
a = 8'd157; b = 8'd36;  #10 
a = 8'd157; b = 8'd37;  #10 
a = 8'd157; b = 8'd38;  #10 
a = 8'd157; b = 8'd39;  #10 
a = 8'd157; b = 8'd40;  #10 
a = 8'd157; b = 8'd41;  #10 
a = 8'd157; b = 8'd42;  #10 
a = 8'd157; b = 8'd43;  #10 
a = 8'd157; b = 8'd44;  #10 
a = 8'd157; b = 8'd45;  #10 
a = 8'd157; b = 8'd46;  #10 
a = 8'd157; b = 8'd47;  #10 
a = 8'd157; b = 8'd48;  #10 
a = 8'd157; b = 8'd49;  #10 
a = 8'd157; b = 8'd50;  #10 
a = 8'd157; b = 8'd51;  #10 
a = 8'd157; b = 8'd52;  #10 
a = 8'd157; b = 8'd53;  #10 
a = 8'd157; b = 8'd54;  #10 
a = 8'd157; b = 8'd55;  #10 
a = 8'd157; b = 8'd56;  #10 
a = 8'd157; b = 8'd57;  #10 
a = 8'd157; b = 8'd58;  #10 
a = 8'd157; b = 8'd59;  #10 
a = 8'd157; b = 8'd60;  #10 
a = 8'd157; b = 8'd61;  #10 
a = 8'd157; b = 8'd62;  #10 
a = 8'd157; b = 8'd63;  #10 
a = 8'd157; b = 8'd64;  #10 
a = 8'd157; b = 8'd65;  #10 
a = 8'd157; b = 8'd66;  #10 
a = 8'd157; b = 8'd67;  #10 
a = 8'd157; b = 8'd68;  #10 
a = 8'd157; b = 8'd69;  #10 
a = 8'd157; b = 8'd70;  #10 
a = 8'd157; b = 8'd71;  #10 
a = 8'd157; b = 8'd72;  #10 
a = 8'd157; b = 8'd73;  #10 
a = 8'd157; b = 8'd74;  #10 
a = 8'd157; b = 8'd75;  #10 
a = 8'd157; b = 8'd76;  #10 
a = 8'd157; b = 8'd77;  #10 
a = 8'd157; b = 8'd78;  #10 
a = 8'd157; b = 8'd79;  #10 
a = 8'd157; b = 8'd80;  #10 
a = 8'd157; b = 8'd81;  #10 
a = 8'd157; b = 8'd82;  #10 
a = 8'd157; b = 8'd83;  #10 
a = 8'd157; b = 8'd84;  #10 
a = 8'd157; b = 8'd85;  #10 
a = 8'd157; b = 8'd86;  #10 
a = 8'd157; b = 8'd87;  #10 
a = 8'd157; b = 8'd88;  #10 
a = 8'd157; b = 8'd89;  #10 
a = 8'd157; b = 8'd90;  #10 
a = 8'd157; b = 8'd91;  #10 
a = 8'd157; b = 8'd92;  #10 
a = 8'd157; b = 8'd93;  #10 
a = 8'd157; b = 8'd94;  #10 
a = 8'd157; b = 8'd95;  #10 
a = 8'd157; b = 8'd96;  #10 
a = 8'd157; b = 8'd97;  #10 
a = 8'd157; b = 8'd98;  #10 
a = 8'd157; b = 8'd99;  #10 
a = 8'd157; b = 8'd100;  #10 
a = 8'd157; b = 8'd101;  #10 
a = 8'd157; b = 8'd102;  #10 
a = 8'd157; b = 8'd103;  #10 
a = 8'd157; b = 8'd104;  #10 
a = 8'd157; b = 8'd105;  #10 
a = 8'd157; b = 8'd106;  #10 
a = 8'd157; b = 8'd107;  #10 
a = 8'd157; b = 8'd108;  #10 
a = 8'd157; b = 8'd109;  #10 
a = 8'd157; b = 8'd110;  #10 
a = 8'd157; b = 8'd111;  #10 
a = 8'd157; b = 8'd112;  #10 
a = 8'd157; b = 8'd113;  #10 
a = 8'd157; b = 8'd114;  #10 
a = 8'd157; b = 8'd115;  #10 
a = 8'd157; b = 8'd116;  #10 
a = 8'd157; b = 8'd117;  #10 
a = 8'd157; b = 8'd118;  #10 
a = 8'd157; b = 8'd119;  #10 
a = 8'd157; b = 8'd120;  #10 
a = 8'd157; b = 8'd121;  #10 
a = 8'd157; b = 8'd122;  #10 
a = 8'd157; b = 8'd123;  #10 
a = 8'd157; b = 8'd124;  #10 
a = 8'd157; b = 8'd125;  #10 
a = 8'd157; b = 8'd126;  #10 
a = 8'd157; b = 8'd127;  #10 
a = 8'd157; b = 8'd128;  #10 
a = 8'd157; b = 8'd129;  #10 
a = 8'd157; b = 8'd130;  #10 
a = 8'd157; b = 8'd131;  #10 
a = 8'd157; b = 8'd132;  #10 
a = 8'd157; b = 8'd133;  #10 
a = 8'd157; b = 8'd134;  #10 
a = 8'd157; b = 8'd135;  #10 
a = 8'd157; b = 8'd136;  #10 
a = 8'd157; b = 8'd137;  #10 
a = 8'd157; b = 8'd138;  #10 
a = 8'd157; b = 8'd139;  #10 
a = 8'd157; b = 8'd140;  #10 
a = 8'd157; b = 8'd141;  #10 
a = 8'd157; b = 8'd142;  #10 
a = 8'd157; b = 8'd143;  #10 
a = 8'd157; b = 8'd144;  #10 
a = 8'd157; b = 8'd145;  #10 
a = 8'd157; b = 8'd146;  #10 
a = 8'd157; b = 8'd147;  #10 
a = 8'd157; b = 8'd148;  #10 
a = 8'd157; b = 8'd149;  #10 
a = 8'd157; b = 8'd150;  #10 
a = 8'd157; b = 8'd151;  #10 
a = 8'd157; b = 8'd152;  #10 
a = 8'd157; b = 8'd153;  #10 
a = 8'd157; b = 8'd154;  #10 
a = 8'd157; b = 8'd155;  #10 
a = 8'd157; b = 8'd156;  #10 
a = 8'd157; b = 8'd157;  #10 
a = 8'd157; b = 8'd158;  #10 
a = 8'd157; b = 8'd159;  #10 
a = 8'd157; b = 8'd160;  #10 
a = 8'd157; b = 8'd161;  #10 
a = 8'd157; b = 8'd162;  #10 
a = 8'd157; b = 8'd163;  #10 
a = 8'd157; b = 8'd164;  #10 
a = 8'd157; b = 8'd165;  #10 
a = 8'd157; b = 8'd166;  #10 
a = 8'd157; b = 8'd167;  #10 
a = 8'd157; b = 8'd168;  #10 
a = 8'd157; b = 8'd169;  #10 
a = 8'd157; b = 8'd170;  #10 
a = 8'd157; b = 8'd171;  #10 
a = 8'd157; b = 8'd172;  #10 
a = 8'd157; b = 8'd173;  #10 
a = 8'd157; b = 8'd174;  #10 
a = 8'd157; b = 8'd175;  #10 
a = 8'd157; b = 8'd176;  #10 
a = 8'd157; b = 8'd177;  #10 
a = 8'd157; b = 8'd178;  #10 
a = 8'd157; b = 8'd179;  #10 
a = 8'd157; b = 8'd180;  #10 
a = 8'd157; b = 8'd181;  #10 
a = 8'd157; b = 8'd182;  #10 
a = 8'd157; b = 8'd183;  #10 
a = 8'd157; b = 8'd184;  #10 
a = 8'd157; b = 8'd185;  #10 
a = 8'd157; b = 8'd186;  #10 
a = 8'd157; b = 8'd187;  #10 
a = 8'd157; b = 8'd188;  #10 
a = 8'd157; b = 8'd189;  #10 
a = 8'd157; b = 8'd190;  #10 
a = 8'd157; b = 8'd191;  #10 
a = 8'd157; b = 8'd192;  #10 
a = 8'd157; b = 8'd193;  #10 
a = 8'd157; b = 8'd194;  #10 
a = 8'd157; b = 8'd195;  #10 
a = 8'd157; b = 8'd196;  #10 
a = 8'd157; b = 8'd197;  #10 
a = 8'd157; b = 8'd198;  #10 
a = 8'd157; b = 8'd199;  #10 
a = 8'd157; b = 8'd200;  #10 
a = 8'd157; b = 8'd201;  #10 
a = 8'd157; b = 8'd202;  #10 
a = 8'd157; b = 8'd203;  #10 
a = 8'd157; b = 8'd204;  #10 
a = 8'd157; b = 8'd205;  #10 
a = 8'd157; b = 8'd206;  #10 
a = 8'd157; b = 8'd207;  #10 
a = 8'd157; b = 8'd208;  #10 
a = 8'd157; b = 8'd209;  #10 
a = 8'd157; b = 8'd210;  #10 
a = 8'd157; b = 8'd211;  #10 
a = 8'd157; b = 8'd212;  #10 
a = 8'd157; b = 8'd213;  #10 
a = 8'd157; b = 8'd214;  #10 
a = 8'd157; b = 8'd215;  #10 
a = 8'd157; b = 8'd216;  #10 
a = 8'd157; b = 8'd217;  #10 
a = 8'd157; b = 8'd218;  #10 
a = 8'd157; b = 8'd219;  #10 
a = 8'd157; b = 8'd220;  #10 
a = 8'd157; b = 8'd221;  #10 
a = 8'd157; b = 8'd222;  #10 
a = 8'd157; b = 8'd223;  #10 
a = 8'd157; b = 8'd224;  #10 
a = 8'd157; b = 8'd225;  #10 
a = 8'd157; b = 8'd226;  #10 
a = 8'd157; b = 8'd227;  #10 
a = 8'd157; b = 8'd228;  #10 
a = 8'd157; b = 8'd229;  #10 
a = 8'd157; b = 8'd230;  #10 
a = 8'd157; b = 8'd231;  #10 
a = 8'd157; b = 8'd232;  #10 
a = 8'd157; b = 8'd233;  #10 
a = 8'd157; b = 8'd234;  #10 
a = 8'd157; b = 8'd235;  #10 
a = 8'd157; b = 8'd236;  #10 
a = 8'd157; b = 8'd237;  #10 
a = 8'd157; b = 8'd238;  #10 
a = 8'd157; b = 8'd239;  #10 
a = 8'd157; b = 8'd240;  #10 
a = 8'd157; b = 8'd241;  #10 
a = 8'd157; b = 8'd242;  #10 
a = 8'd157; b = 8'd243;  #10 
a = 8'd157; b = 8'd244;  #10 
a = 8'd157; b = 8'd245;  #10 
a = 8'd157; b = 8'd246;  #10 
a = 8'd157; b = 8'd247;  #10 
a = 8'd157; b = 8'd248;  #10 
a = 8'd157; b = 8'd249;  #10 
a = 8'd157; b = 8'd250;  #10 
a = 8'd157; b = 8'd251;  #10 
a = 8'd157; b = 8'd252;  #10 
a = 8'd157; b = 8'd253;  #10 
a = 8'd157; b = 8'd254;  #10 
a = 8'd157; b = 8'd255;  #10 
a = 8'd158; b = 8'd0;  #10 
a = 8'd158; b = 8'd1;  #10 
a = 8'd158; b = 8'd2;  #10 
a = 8'd158; b = 8'd3;  #10 
a = 8'd158; b = 8'd4;  #10 
a = 8'd158; b = 8'd5;  #10 
a = 8'd158; b = 8'd6;  #10 
a = 8'd158; b = 8'd7;  #10 
a = 8'd158; b = 8'd8;  #10 
a = 8'd158; b = 8'd9;  #10 
a = 8'd158; b = 8'd10;  #10 
a = 8'd158; b = 8'd11;  #10 
a = 8'd158; b = 8'd12;  #10 
a = 8'd158; b = 8'd13;  #10 
a = 8'd158; b = 8'd14;  #10 
a = 8'd158; b = 8'd15;  #10 
a = 8'd158; b = 8'd16;  #10 
a = 8'd158; b = 8'd17;  #10 
a = 8'd158; b = 8'd18;  #10 
a = 8'd158; b = 8'd19;  #10 
a = 8'd158; b = 8'd20;  #10 
a = 8'd158; b = 8'd21;  #10 
a = 8'd158; b = 8'd22;  #10 
a = 8'd158; b = 8'd23;  #10 
a = 8'd158; b = 8'd24;  #10 
a = 8'd158; b = 8'd25;  #10 
a = 8'd158; b = 8'd26;  #10 
a = 8'd158; b = 8'd27;  #10 
a = 8'd158; b = 8'd28;  #10 
a = 8'd158; b = 8'd29;  #10 
a = 8'd158; b = 8'd30;  #10 
a = 8'd158; b = 8'd31;  #10 
a = 8'd158; b = 8'd32;  #10 
a = 8'd158; b = 8'd33;  #10 
a = 8'd158; b = 8'd34;  #10 
a = 8'd158; b = 8'd35;  #10 
a = 8'd158; b = 8'd36;  #10 
a = 8'd158; b = 8'd37;  #10 
a = 8'd158; b = 8'd38;  #10 
a = 8'd158; b = 8'd39;  #10 
a = 8'd158; b = 8'd40;  #10 
a = 8'd158; b = 8'd41;  #10 
a = 8'd158; b = 8'd42;  #10 
a = 8'd158; b = 8'd43;  #10 
a = 8'd158; b = 8'd44;  #10 
a = 8'd158; b = 8'd45;  #10 
a = 8'd158; b = 8'd46;  #10 
a = 8'd158; b = 8'd47;  #10 
a = 8'd158; b = 8'd48;  #10 
a = 8'd158; b = 8'd49;  #10 
a = 8'd158; b = 8'd50;  #10 
a = 8'd158; b = 8'd51;  #10 
a = 8'd158; b = 8'd52;  #10 
a = 8'd158; b = 8'd53;  #10 
a = 8'd158; b = 8'd54;  #10 
a = 8'd158; b = 8'd55;  #10 
a = 8'd158; b = 8'd56;  #10 
a = 8'd158; b = 8'd57;  #10 
a = 8'd158; b = 8'd58;  #10 
a = 8'd158; b = 8'd59;  #10 
a = 8'd158; b = 8'd60;  #10 
a = 8'd158; b = 8'd61;  #10 
a = 8'd158; b = 8'd62;  #10 
a = 8'd158; b = 8'd63;  #10 
a = 8'd158; b = 8'd64;  #10 
a = 8'd158; b = 8'd65;  #10 
a = 8'd158; b = 8'd66;  #10 
a = 8'd158; b = 8'd67;  #10 
a = 8'd158; b = 8'd68;  #10 
a = 8'd158; b = 8'd69;  #10 
a = 8'd158; b = 8'd70;  #10 
a = 8'd158; b = 8'd71;  #10 
a = 8'd158; b = 8'd72;  #10 
a = 8'd158; b = 8'd73;  #10 
a = 8'd158; b = 8'd74;  #10 
a = 8'd158; b = 8'd75;  #10 
a = 8'd158; b = 8'd76;  #10 
a = 8'd158; b = 8'd77;  #10 
a = 8'd158; b = 8'd78;  #10 
a = 8'd158; b = 8'd79;  #10 
a = 8'd158; b = 8'd80;  #10 
a = 8'd158; b = 8'd81;  #10 
a = 8'd158; b = 8'd82;  #10 
a = 8'd158; b = 8'd83;  #10 
a = 8'd158; b = 8'd84;  #10 
a = 8'd158; b = 8'd85;  #10 
a = 8'd158; b = 8'd86;  #10 
a = 8'd158; b = 8'd87;  #10 
a = 8'd158; b = 8'd88;  #10 
a = 8'd158; b = 8'd89;  #10 
a = 8'd158; b = 8'd90;  #10 
a = 8'd158; b = 8'd91;  #10 
a = 8'd158; b = 8'd92;  #10 
a = 8'd158; b = 8'd93;  #10 
a = 8'd158; b = 8'd94;  #10 
a = 8'd158; b = 8'd95;  #10 
a = 8'd158; b = 8'd96;  #10 
a = 8'd158; b = 8'd97;  #10 
a = 8'd158; b = 8'd98;  #10 
a = 8'd158; b = 8'd99;  #10 
a = 8'd158; b = 8'd100;  #10 
a = 8'd158; b = 8'd101;  #10 
a = 8'd158; b = 8'd102;  #10 
a = 8'd158; b = 8'd103;  #10 
a = 8'd158; b = 8'd104;  #10 
a = 8'd158; b = 8'd105;  #10 
a = 8'd158; b = 8'd106;  #10 
a = 8'd158; b = 8'd107;  #10 
a = 8'd158; b = 8'd108;  #10 
a = 8'd158; b = 8'd109;  #10 
a = 8'd158; b = 8'd110;  #10 
a = 8'd158; b = 8'd111;  #10 
a = 8'd158; b = 8'd112;  #10 
a = 8'd158; b = 8'd113;  #10 
a = 8'd158; b = 8'd114;  #10 
a = 8'd158; b = 8'd115;  #10 
a = 8'd158; b = 8'd116;  #10 
a = 8'd158; b = 8'd117;  #10 
a = 8'd158; b = 8'd118;  #10 
a = 8'd158; b = 8'd119;  #10 
a = 8'd158; b = 8'd120;  #10 
a = 8'd158; b = 8'd121;  #10 
a = 8'd158; b = 8'd122;  #10 
a = 8'd158; b = 8'd123;  #10 
a = 8'd158; b = 8'd124;  #10 
a = 8'd158; b = 8'd125;  #10 
a = 8'd158; b = 8'd126;  #10 
a = 8'd158; b = 8'd127;  #10 
a = 8'd158; b = 8'd128;  #10 
a = 8'd158; b = 8'd129;  #10 
a = 8'd158; b = 8'd130;  #10 
a = 8'd158; b = 8'd131;  #10 
a = 8'd158; b = 8'd132;  #10 
a = 8'd158; b = 8'd133;  #10 
a = 8'd158; b = 8'd134;  #10 
a = 8'd158; b = 8'd135;  #10 
a = 8'd158; b = 8'd136;  #10 
a = 8'd158; b = 8'd137;  #10 
a = 8'd158; b = 8'd138;  #10 
a = 8'd158; b = 8'd139;  #10 
a = 8'd158; b = 8'd140;  #10 
a = 8'd158; b = 8'd141;  #10 
a = 8'd158; b = 8'd142;  #10 
a = 8'd158; b = 8'd143;  #10 
a = 8'd158; b = 8'd144;  #10 
a = 8'd158; b = 8'd145;  #10 
a = 8'd158; b = 8'd146;  #10 
a = 8'd158; b = 8'd147;  #10 
a = 8'd158; b = 8'd148;  #10 
a = 8'd158; b = 8'd149;  #10 
a = 8'd158; b = 8'd150;  #10 
a = 8'd158; b = 8'd151;  #10 
a = 8'd158; b = 8'd152;  #10 
a = 8'd158; b = 8'd153;  #10 
a = 8'd158; b = 8'd154;  #10 
a = 8'd158; b = 8'd155;  #10 
a = 8'd158; b = 8'd156;  #10 
a = 8'd158; b = 8'd157;  #10 
a = 8'd158; b = 8'd158;  #10 
a = 8'd158; b = 8'd159;  #10 
a = 8'd158; b = 8'd160;  #10 
a = 8'd158; b = 8'd161;  #10 
a = 8'd158; b = 8'd162;  #10 
a = 8'd158; b = 8'd163;  #10 
a = 8'd158; b = 8'd164;  #10 
a = 8'd158; b = 8'd165;  #10 
a = 8'd158; b = 8'd166;  #10 
a = 8'd158; b = 8'd167;  #10 
a = 8'd158; b = 8'd168;  #10 
a = 8'd158; b = 8'd169;  #10 
a = 8'd158; b = 8'd170;  #10 
a = 8'd158; b = 8'd171;  #10 
a = 8'd158; b = 8'd172;  #10 
a = 8'd158; b = 8'd173;  #10 
a = 8'd158; b = 8'd174;  #10 
a = 8'd158; b = 8'd175;  #10 
a = 8'd158; b = 8'd176;  #10 
a = 8'd158; b = 8'd177;  #10 
a = 8'd158; b = 8'd178;  #10 
a = 8'd158; b = 8'd179;  #10 
a = 8'd158; b = 8'd180;  #10 
a = 8'd158; b = 8'd181;  #10 
a = 8'd158; b = 8'd182;  #10 
a = 8'd158; b = 8'd183;  #10 
a = 8'd158; b = 8'd184;  #10 
a = 8'd158; b = 8'd185;  #10 
a = 8'd158; b = 8'd186;  #10 
a = 8'd158; b = 8'd187;  #10 
a = 8'd158; b = 8'd188;  #10 
a = 8'd158; b = 8'd189;  #10 
a = 8'd158; b = 8'd190;  #10 
a = 8'd158; b = 8'd191;  #10 
a = 8'd158; b = 8'd192;  #10 
a = 8'd158; b = 8'd193;  #10 
a = 8'd158; b = 8'd194;  #10 
a = 8'd158; b = 8'd195;  #10 
a = 8'd158; b = 8'd196;  #10 
a = 8'd158; b = 8'd197;  #10 
a = 8'd158; b = 8'd198;  #10 
a = 8'd158; b = 8'd199;  #10 
a = 8'd158; b = 8'd200;  #10 
a = 8'd158; b = 8'd201;  #10 
a = 8'd158; b = 8'd202;  #10 
a = 8'd158; b = 8'd203;  #10 
a = 8'd158; b = 8'd204;  #10 
a = 8'd158; b = 8'd205;  #10 
a = 8'd158; b = 8'd206;  #10 
a = 8'd158; b = 8'd207;  #10 
a = 8'd158; b = 8'd208;  #10 
a = 8'd158; b = 8'd209;  #10 
a = 8'd158; b = 8'd210;  #10 
a = 8'd158; b = 8'd211;  #10 
a = 8'd158; b = 8'd212;  #10 
a = 8'd158; b = 8'd213;  #10 
a = 8'd158; b = 8'd214;  #10 
a = 8'd158; b = 8'd215;  #10 
a = 8'd158; b = 8'd216;  #10 
a = 8'd158; b = 8'd217;  #10 
a = 8'd158; b = 8'd218;  #10 
a = 8'd158; b = 8'd219;  #10 
a = 8'd158; b = 8'd220;  #10 
a = 8'd158; b = 8'd221;  #10 
a = 8'd158; b = 8'd222;  #10 
a = 8'd158; b = 8'd223;  #10 
a = 8'd158; b = 8'd224;  #10 
a = 8'd158; b = 8'd225;  #10 
a = 8'd158; b = 8'd226;  #10 
a = 8'd158; b = 8'd227;  #10 
a = 8'd158; b = 8'd228;  #10 
a = 8'd158; b = 8'd229;  #10 
a = 8'd158; b = 8'd230;  #10 
a = 8'd158; b = 8'd231;  #10 
a = 8'd158; b = 8'd232;  #10 
a = 8'd158; b = 8'd233;  #10 
a = 8'd158; b = 8'd234;  #10 
a = 8'd158; b = 8'd235;  #10 
a = 8'd158; b = 8'd236;  #10 
a = 8'd158; b = 8'd237;  #10 
a = 8'd158; b = 8'd238;  #10 
a = 8'd158; b = 8'd239;  #10 
a = 8'd158; b = 8'd240;  #10 
a = 8'd158; b = 8'd241;  #10 
a = 8'd158; b = 8'd242;  #10 
a = 8'd158; b = 8'd243;  #10 
a = 8'd158; b = 8'd244;  #10 
a = 8'd158; b = 8'd245;  #10 
a = 8'd158; b = 8'd246;  #10 
a = 8'd158; b = 8'd247;  #10 
a = 8'd158; b = 8'd248;  #10 
a = 8'd158; b = 8'd249;  #10 
a = 8'd158; b = 8'd250;  #10 
a = 8'd158; b = 8'd251;  #10 
a = 8'd158; b = 8'd252;  #10 
a = 8'd158; b = 8'd253;  #10 
a = 8'd158; b = 8'd254;  #10 
a = 8'd158; b = 8'd255;  #10 
a = 8'd159; b = 8'd0;  #10 
a = 8'd159; b = 8'd1;  #10 
a = 8'd159; b = 8'd2;  #10 
a = 8'd159; b = 8'd3;  #10 
a = 8'd159; b = 8'd4;  #10 
a = 8'd159; b = 8'd5;  #10 
a = 8'd159; b = 8'd6;  #10 
a = 8'd159; b = 8'd7;  #10 
a = 8'd159; b = 8'd8;  #10 
a = 8'd159; b = 8'd9;  #10 
a = 8'd159; b = 8'd10;  #10 
a = 8'd159; b = 8'd11;  #10 
a = 8'd159; b = 8'd12;  #10 
a = 8'd159; b = 8'd13;  #10 
a = 8'd159; b = 8'd14;  #10 
a = 8'd159; b = 8'd15;  #10 
a = 8'd159; b = 8'd16;  #10 
a = 8'd159; b = 8'd17;  #10 
a = 8'd159; b = 8'd18;  #10 
a = 8'd159; b = 8'd19;  #10 
a = 8'd159; b = 8'd20;  #10 
a = 8'd159; b = 8'd21;  #10 
a = 8'd159; b = 8'd22;  #10 
a = 8'd159; b = 8'd23;  #10 
a = 8'd159; b = 8'd24;  #10 
a = 8'd159; b = 8'd25;  #10 
a = 8'd159; b = 8'd26;  #10 
a = 8'd159; b = 8'd27;  #10 
a = 8'd159; b = 8'd28;  #10 
a = 8'd159; b = 8'd29;  #10 
a = 8'd159; b = 8'd30;  #10 
a = 8'd159; b = 8'd31;  #10 
a = 8'd159; b = 8'd32;  #10 
a = 8'd159; b = 8'd33;  #10 
a = 8'd159; b = 8'd34;  #10 
a = 8'd159; b = 8'd35;  #10 
a = 8'd159; b = 8'd36;  #10 
a = 8'd159; b = 8'd37;  #10 
a = 8'd159; b = 8'd38;  #10 
a = 8'd159; b = 8'd39;  #10 
a = 8'd159; b = 8'd40;  #10 
a = 8'd159; b = 8'd41;  #10 
a = 8'd159; b = 8'd42;  #10 
a = 8'd159; b = 8'd43;  #10 
a = 8'd159; b = 8'd44;  #10 
a = 8'd159; b = 8'd45;  #10 
a = 8'd159; b = 8'd46;  #10 
a = 8'd159; b = 8'd47;  #10 
a = 8'd159; b = 8'd48;  #10 
a = 8'd159; b = 8'd49;  #10 
a = 8'd159; b = 8'd50;  #10 
a = 8'd159; b = 8'd51;  #10 
a = 8'd159; b = 8'd52;  #10 
a = 8'd159; b = 8'd53;  #10 
a = 8'd159; b = 8'd54;  #10 
a = 8'd159; b = 8'd55;  #10 
a = 8'd159; b = 8'd56;  #10 
a = 8'd159; b = 8'd57;  #10 
a = 8'd159; b = 8'd58;  #10 
a = 8'd159; b = 8'd59;  #10 
a = 8'd159; b = 8'd60;  #10 
a = 8'd159; b = 8'd61;  #10 
a = 8'd159; b = 8'd62;  #10 
a = 8'd159; b = 8'd63;  #10 
a = 8'd159; b = 8'd64;  #10 
a = 8'd159; b = 8'd65;  #10 
a = 8'd159; b = 8'd66;  #10 
a = 8'd159; b = 8'd67;  #10 
a = 8'd159; b = 8'd68;  #10 
a = 8'd159; b = 8'd69;  #10 
a = 8'd159; b = 8'd70;  #10 
a = 8'd159; b = 8'd71;  #10 
a = 8'd159; b = 8'd72;  #10 
a = 8'd159; b = 8'd73;  #10 
a = 8'd159; b = 8'd74;  #10 
a = 8'd159; b = 8'd75;  #10 
a = 8'd159; b = 8'd76;  #10 
a = 8'd159; b = 8'd77;  #10 
a = 8'd159; b = 8'd78;  #10 
a = 8'd159; b = 8'd79;  #10 
a = 8'd159; b = 8'd80;  #10 
a = 8'd159; b = 8'd81;  #10 
a = 8'd159; b = 8'd82;  #10 
a = 8'd159; b = 8'd83;  #10 
a = 8'd159; b = 8'd84;  #10 
a = 8'd159; b = 8'd85;  #10 
a = 8'd159; b = 8'd86;  #10 
a = 8'd159; b = 8'd87;  #10 
a = 8'd159; b = 8'd88;  #10 
a = 8'd159; b = 8'd89;  #10 
a = 8'd159; b = 8'd90;  #10 
a = 8'd159; b = 8'd91;  #10 
a = 8'd159; b = 8'd92;  #10 
a = 8'd159; b = 8'd93;  #10 
a = 8'd159; b = 8'd94;  #10 
a = 8'd159; b = 8'd95;  #10 
a = 8'd159; b = 8'd96;  #10 
a = 8'd159; b = 8'd97;  #10 
a = 8'd159; b = 8'd98;  #10 
a = 8'd159; b = 8'd99;  #10 
a = 8'd159; b = 8'd100;  #10 
a = 8'd159; b = 8'd101;  #10 
a = 8'd159; b = 8'd102;  #10 
a = 8'd159; b = 8'd103;  #10 
a = 8'd159; b = 8'd104;  #10 
a = 8'd159; b = 8'd105;  #10 
a = 8'd159; b = 8'd106;  #10 
a = 8'd159; b = 8'd107;  #10 
a = 8'd159; b = 8'd108;  #10 
a = 8'd159; b = 8'd109;  #10 
a = 8'd159; b = 8'd110;  #10 
a = 8'd159; b = 8'd111;  #10 
a = 8'd159; b = 8'd112;  #10 
a = 8'd159; b = 8'd113;  #10 
a = 8'd159; b = 8'd114;  #10 
a = 8'd159; b = 8'd115;  #10 
a = 8'd159; b = 8'd116;  #10 
a = 8'd159; b = 8'd117;  #10 
a = 8'd159; b = 8'd118;  #10 
a = 8'd159; b = 8'd119;  #10 
a = 8'd159; b = 8'd120;  #10 
a = 8'd159; b = 8'd121;  #10 
a = 8'd159; b = 8'd122;  #10 
a = 8'd159; b = 8'd123;  #10 
a = 8'd159; b = 8'd124;  #10 
a = 8'd159; b = 8'd125;  #10 
a = 8'd159; b = 8'd126;  #10 
a = 8'd159; b = 8'd127;  #10 
a = 8'd159; b = 8'd128;  #10 
a = 8'd159; b = 8'd129;  #10 
a = 8'd159; b = 8'd130;  #10 
a = 8'd159; b = 8'd131;  #10 
a = 8'd159; b = 8'd132;  #10 
a = 8'd159; b = 8'd133;  #10 
a = 8'd159; b = 8'd134;  #10 
a = 8'd159; b = 8'd135;  #10 
a = 8'd159; b = 8'd136;  #10 
a = 8'd159; b = 8'd137;  #10 
a = 8'd159; b = 8'd138;  #10 
a = 8'd159; b = 8'd139;  #10 
a = 8'd159; b = 8'd140;  #10 
a = 8'd159; b = 8'd141;  #10 
a = 8'd159; b = 8'd142;  #10 
a = 8'd159; b = 8'd143;  #10 
a = 8'd159; b = 8'd144;  #10 
a = 8'd159; b = 8'd145;  #10 
a = 8'd159; b = 8'd146;  #10 
a = 8'd159; b = 8'd147;  #10 
a = 8'd159; b = 8'd148;  #10 
a = 8'd159; b = 8'd149;  #10 
a = 8'd159; b = 8'd150;  #10 
a = 8'd159; b = 8'd151;  #10 
a = 8'd159; b = 8'd152;  #10 
a = 8'd159; b = 8'd153;  #10 
a = 8'd159; b = 8'd154;  #10 
a = 8'd159; b = 8'd155;  #10 
a = 8'd159; b = 8'd156;  #10 
a = 8'd159; b = 8'd157;  #10 
a = 8'd159; b = 8'd158;  #10 
a = 8'd159; b = 8'd159;  #10 
a = 8'd159; b = 8'd160;  #10 
a = 8'd159; b = 8'd161;  #10 
a = 8'd159; b = 8'd162;  #10 
a = 8'd159; b = 8'd163;  #10 
a = 8'd159; b = 8'd164;  #10 
a = 8'd159; b = 8'd165;  #10 
a = 8'd159; b = 8'd166;  #10 
a = 8'd159; b = 8'd167;  #10 
a = 8'd159; b = 8'd168;  #10 
a = 8'd159; b = 8'd169;  #10 
a = 8'd159; b = 8'd170;  #10 
a = 8'd159; b = 8'd171;  #10 
a = 8'd159; b = 8'd172;  #10 
a = 8'd159; b = 8'd173;  #10 
a = 8'd159; b = 8'd174;  #10 
a = 8'd159; b = 8'd175;  #10 
a = 8'd159; b = 8'd176;  #10 
a = 8'd159; b = 8'd177;  #10 
a = 8'd159; b = 8'd178;  #10 
a = 8'd159; b = 8'd179;  #10 
a = 8'd159; b = 8'd180;  #10 
a = 8'd159; b = 8'd181;  #10 
a = 8'd159; b = 8'd182;  #10 
a = 8'd159; b = 8'd183;  #10 
a = 8'd159; b = 8'd184;  #10 
a = 8'd159; b = 8'd185;  #10 
a = 8'd159; b = 8'd186;  #10 
a = 8'd159; b = 8'd187;  #10 
a = 8'd159; b = 8'd188;  #10 
a = 8'd159; b = 8'd189;  #10 
a = 8'd159; b = 8'd190;  #10 
a = 8'd159; b = 8'd191;  #10 
a = 8'd159; b = 8'd192;  #10 
a = 8'd159; b = 8'd193;  #10 
a = 8'd159; b = 8'd194;  #10 
a = 8'd159; b = 8'd195;  #10 
a = 8'd159; b = 8'd196;  #10 
a = 8'd159; b = 8'd197;  #10 
a = 8'd159; b = 8'd198;  #10 
a = 8'd159; b = 8'd199;  #10 
a = 8'd159; b = 8'd200;  #10 
a = 8'd159; b = 8'd201;  #10 
a = 8'd159; b = 8'd202;  #10 
a = 8'd159; b = 8'd203;  #10 
a = 8'd159; b = 8'd204;  #10 
a = 8'd159; b = 8'd205;  #10 
a = 8'd159; b = 8'd206;  #10 
a = 8'd159; b = 8'd207;  #10 
a = 8'd159; b = 8'd208;  #10 
a = 8'd159; b = 8'd209;  #10 
a = 8'd159; b = 8'd210;  #10 
a = 8'd159; b = 8'd211;  #10 
a = 8'd159; b = 8'd212;  #10 
a = 8'd159; b = 8'd213;  #10 
a = 8'd159; b = 8'd214;  #10 
a = 8'd159; b = 8'd215;  #10 
a = 8'd159; b = 8'd216;  #10 
a = 8'd159; b = 8'd217;  #10 
a = 8'd159; b = 8'd218;  #10 
a = 8'd159; b = 8'd219;  #10 
a = 8'd159; b = 8'd220;  #10 
a = 8'd159; b = 8'd221;  #10 
a = 8'd159; b = 8'd222;  #10 
a = 8'd159; b = 8'd223;  #10 
a = 8'd159; b = 8'd224;  #10 
a = 8'd159; b = 8'd225;  #10 
a = 8'd159; b = 8'd226;  #10 
a = 8'd159; b = 8'd227;  #10 
a = 8'd159; b = 8'd228;  #10 
a = 8'd159; b = 8'd229;  #10 
a = 8'd159; b = 8'd230;  #10 
a = 8'd159; b = 8'd231;  #10 
a = 8'd159; b = 8'd232;  #10 
a = 8'd159; b = 8'd233;  #10 
a = 8'd159; b = 8'd234;  #10 
a = 8'd159; b = 8'd235;  #10 
a = 8'd159; b = 8'd236;  #10 
a = 8'd159; b = 8'd237;  #10 
a = 8'd159; b = 8'd238;  #10 
a = 8'd159; b = 8'd239;  #10 
a = 8'd159; b = 8'd240;  #10 
a = 8'd159; b = 8'd241;  #10 
a = 8'd159; b = 8'd242;  #10 
a = 8'd159; b = 8'd243;  #10 
a = 8'd159; b = 8'd244;  #10 
a = 8'd159; b = 8'd245;  #10 
a = 8'd159; b = 8'd246;  #10 
a = 8'd159; b = 8'd247;  #10 
a = 8'd159; b = 8'd248;  #10 
a = 8'd159; b = 8'd249;  #10 
a = 8'd159; b = 8'd250;  #10 
a = 8'd159; b = 8'd251;  #10 
a = 8'd159; b = 8'd252;  #10 
a = 8'd159; b = 8'd253;  #10 
a = 8'd159; b = 8'd254;  #10 
a = 8'd159; b = 8'd255;  #10 
a = 8'd160; b = 8'd0;  #10 
a = 8'd160; b = 8'd1;  #10 
a = 8'd160; b = 8'd2;  #10 
a = 8'd160; b = 8'd3;  #10 
a = 8'd160; b = 8'd4;  #10 
a = 8'd160; b = 8'd5;  #10 
a = 8'd160; b = 8'd6;  #10 
a = 8'd160; b = 8'd7;  #10 
a = 8'd160; b = 8'd8;  #10 
a = 8'd160; b = 8'd9;  #10 
a = 8'd160; b = 8'd10;  #10 
a = 8'd160; b = 8'd11;  #10 
a = 8'd160; b = 8'd12;  #10 
a = 8'd160; b = 8'd13;  #10 
a = 8'd160; b = 8'd14;  #10 
a = 8'd160; b = 8'd15;  #10 
a = 8'd160; b = 8'd16;  #10 
a = 8'd160; b = 8'd17;  #10 
a = 8'd160; b = 8'd18;  #10 
a = 8'd160; b = 8'd19;  #10 
a = 8'd160; b = 8'd20;  #10 
a = 8'd160; b = 8'd21;  #10 
a = 8'd160; b = 8'd22;  #10 
a = 8'd160; b = 8'd23;  #10 
a = 8'd160; b = 8'd24;  #10 
a = 8'd160; b = 8'd25;  #10 
a = 8'd160; b = 8'd26;  #10 
a = 8'd160; b = 8'd27;  #10 
a = 8'd160; b = 8'd28;  #10 
a = 8'd160; b = 8'd29;  #10 
a = 8'd160; b = 8'd30;  #10 
a = 8'd160; b = 8'd31;  #10 
a = 8'd160; b = 8'd32;  #10 
a = 8'd160; b = 8'd33;  #10 
a = 8'd160; b = 8'd34;  #10 
a = 8'd160; b = 8'd35;  #10 
a = 8'd160; b = 8'd36;  #10 
a = 8'd160; b = 8'd37;  #10 
a = 8'd160; b = 8'd38;  #10 
a = 8'd160; b = 8'd39;  #10 
a = 8'd160; b = 8'd40;  #10 
a = 8'd160; b = 8'd41;  #10 
a = 8'd160; b = 8'd42;  #10 
a = 8'd160; b = 8'd43;  #10 
a = 8'd160; b = 8'd44;  #10 
a = 8'd160; b = 8'd45;  #10 
a = 8'd160; b = 8'd46;  #10 
a = 8'd160; b = 8'd47;  #10 
a = 8'd160; b = 8'd48;  #10 
a = 8'd160; b = 8'd49;  #10 
a = 8'd160; b = 8'd50;  #10 
a = 8'd160; b = 8'd51;  #10 
a = 8'd160; b = 8'd52;  #10 
a = 8'd160; b = 8'd53;  #10 
a = 8'd160; b = 8'd54;  #10 
a = 8'd160; b = 8'd55;  #10 
a = 8'd160; b = 8'd56;  #10 
a = 8'd160; b = 8'd57;  #10 
a = 8'd160; b = 8'd58;  #10 
a = 8'd160; b = 8'd59;  #10 
a = 8'd160; b = 8'd60;  #10 
a = 8'd160; b = 8'd61;  #10 
a = 8'd160; b = 8'd62;  #10 
a = 8'd160; b = 8'd63;  #10 
a = 8'd160; b = 8'd64;  #10 
a = 8'd160; b = 8'd65;  #10 
a = 8'd160; b = 8'd66;  #10 
a = 8'd160; b = 8'd67;  #10 
a = 8'd160; b = 8'd68;  #10 
a = 8'd160; b = 8'd69;  #10 
a = 8'd160; b = 8'd70;  #10 
a = 8'd160; b = 8'd71;  #10 
a = 8'd160; b = 8'd72;  #10 
a = 8'd160; b = 8'd73;  #10 
a = 8'd160; b = 8'd74;  #10 
a = 8'd160; b = 8'd75;  #10 
a = 8'd160; b = 8'd76;  #10 
a = 8'd160; b = 8'd77;  #10 
a = 8'd160; b = 8'd78;  #10 
a = 8'd160; b = 8'd79;  #10 
a = 8'd160; b = 8'd80;  #10 
a = 8'd160; b = 8'd81;  #10 
a = 8'd160; b = 8'd82;  #10 
a = 8'd160; b = 8'd83;  #10 
a = 8'd160; b = 8'd84;  #10 
a = 8'd160; b = 8'd85;  #10 
a = 8'd160; b = 8'd86;  #10 
a = 8'd160; b = 8'd87;  #10 
a = 8'd160; b = 8'd88;  #10 
a = 8'd160; b = 8'd89;  #10 
a = 8'd160; b = 8'd90;  #10 
a = 8'd160; b = 8'd91;  #10 
a = 8'd160; b = 8'd92;  #10 
a = 8'd160; b = 8'd93;  #10 
a = 8'd160; b = 8'd94;  #10 
a = 8'd160; b = 8'd95;  #10 
a = 8'd160; b = 8'd96;  #10 
a = 8'd160; b = 8'd97;  #10 
a = 8'd160; b = 8'd98;  #10 
a = 8'd160; b = 8'd99;  #10 
a = 8'd160; b = 8'd100;  #10 
a = 8'd160; b = 8'd101;  #10 
a = 8'd160; b = 8'd102;  #10 
a = 8'd160; b = 8'd103;  #10 
a = 8'd160; b = 8'd104;  #10 
a = 8'd160; b = 8'd105;  #10 
a = 8'd160; b = 8'd106;  #10 
a = 8'd160; b = 8'd107;  #10 
a = 8'd160; b = 8'd108;  #10 
a = 8'd160; b = 8'd109;  #10 
a = 8'd160; b = 8'd110;  #10 
a = 8'd160; b = 8'd111;  #10 
a = 8'd160; b = 8'd112;  #10 
a = 8'd160; b = 8'd113;  #10 
a = 8'd160; b = 8'd114;  #10 
a = 8'd160; b = 8'd115;  #10 
a = 8'd160; b = 8'd116;  #10 
a = 8'd160; b = 8'd117;  #10 
a = 8'd160; b = 8'd118;  #10 
a = 8'd160; b = 8'd119;  #10 
a = 8'd160; b = 8'd120;  #10 
a = 8'd160; b = 8'd121;  #10 
a = 8'd160; b = 8'd122;  #10 
a = 8'd160; b = 8'd123;  #10 
a = 8'd160; b = 8'd124;  #10 
a = 8'd160; b = 8'd125;  #10 
a = 8'd160; b = 8'd126;  #10 
a = 8'd160; b = 8'd127;  #10 
a = 8'd160; b = 8'd128;  #10 
a = 8'd160; b = 8'd129;  #10 
a = 8'd160; b = 8'd130;  #10 
a = 8'd160; b = 8'd131;  #10 
a = 8'd160; b = 8'd132;  #10 
a = 8'd160; b = 8'd133;  #10 
a = 8'd160; b = 8'd134;  #10 
a = 8'd160; b = 8'd135;  #10 
a = 8'd160; b = 8'd136;  #10 
a = 8'd160; b = 8'd137;  #10 
a = 8'd160; b = 8'd138;  #10 
a = 8'd160; b = 8'd139;  #10 
a = 8'd160; b = 8'd140;  #10 
a = 8'd160; b = 8'd141;  #10 
a = 8'd160; b = 8'd142;  #10 
a = 8'd160; b = 8'd143;  #10 
a = 8'd160; b = 8'd144;  #10 
a = 8'd160; b = 8'd145;  #10 
a = 8'd160; b = 8'd146;  #10 
a = 8'd160; b = 8'd147;  #10 
a = 8'd160; b = 8'd148;  #10 
a = 8'd160; b = 8'd149;  #10 
a = 8'd160; b = 8'd150;  #10 
a = 8'd160; b = 8'd151;  #10 
a = 8'd160; b = 8'd152;  #10 
a = 8'd160; b = 8'd153;  #10 
a = 8'd160; b = 8'd154;  #10 
a = 8'd160; b = 8'd155;  #10 
a = 8'd160; b = 8'd156;  #10 
a = 8'd160; b = 8'd157;  #10 
a = 8'd160; b = 8'd158;  #10 
a = 8'd160; b = 8'd159;  #10 
a = 8'd160; b = 8'd160;  #10 
a = 8'd160; b = 8'd161;  #10 
a = 8'd160; b = 8'd162;  #10 
a = 8'd160; b = 8'd163;  #10 
a = 8'd160; b = 8'd164;  #10 
a = 8'd160; b = 8'd165;  #10 
a = 8'd160; b = 8'd166;  #10 
a = 8'd160; b = 8'd167;  #10 
a = 8'd160; b = 8'd168;  #10 
a = 8'd160; b = 8'd169;  #10 
a = 8'd160; b = 8'd170;  #10 
a = 8'd160; b = 8'd171;  #10 
a = 8'd160; b = 8'd172;  #10 
a = 8'd160; b = 8'd173;  #10 
a = 8'd160; b = 8'd174;  #10 
a = 8'd160; b = 8'd175;  #10 
a = 8'd160; b = 8'd176;  #10 
a = 8'd160; b = 8'd177;  #10 
a = 8'd160; b = 8'd178;  #10 
a = 8'd160; b = 8'd179;  #10 
a = 8'd160; b = 8'd180;  #10 
a = 8'd160; b = 8'd181;  #10 
a = 8'd160; b = 8'd182;  #10 
a = 8'd160; b = 8'd183;  #10 
a = 8'd160; b = 8'd184;  #10 
a = 8'd160; b = 8'd185;  #10 
a = 8'd160; b = 8'd186;  #10 
a = 8'd160; b = 8'd187;  #10 
a = 8'd160; b = 8'd188;  #10 
a = 8'd160; b = 8'd189;  #10 
a = 8'd160; b = 8'd190;  #10 
a = 8'd160; b = 8'd191;  #10 
a = 8'd160; b = 8'd192;  #10 
a = 8'd160; b = 8'd193;  #10 
a = 8'd160; b = 8'd194;  #10 
a = 8'd160; b = 8'd195;  #10 
a = 8'd160; b = 8'd196;  #10 
a = 8'd160; b = 8'd197;  #10 
a = 8'd160; b = 8'd198;  #10 
a = 8'd160; b = 8'd199;  #10 
a = 8'd160; b = 8'd200;  #10 
a = 8'd160; b = 8'd201;  #10 
a = 8'd160; b = 8'd202;  #10 
a = 8'd160; b = 8'd203;  #10 
a = 8'd160; b = 8'd204;  #10 
a = 8'd160; b = 8'd205;  #10 
a = 8'd160; b = 8'd206;  #10 
a = 8'd160; b = 8'd207;  #10 
a = 8'd160; b = 8'd208;  #10 
a = 8'd160; b = 8'd209;  #10 
a = 8'd160; b = 8'd210;  #10 
a = 8'd160; b = 8'd211;  #10 
a = 8'd160; b = 8'd212;  #10 
a = 8'd160; b = 8'd213;  #10 
a = 8'd160; b = 8'd214;  #10 
a = 8'd160; b = 8'd215;  #10 
a = 8'd160; b = 8'd216;  #10 
a = 8'd160; b = 8'd217;  #10 
a = 8'd160; b = 8'd218;  #10 
a = 8'd160; b = 8'd219;  #10 
a = 8'd160; b = 8'd220;  #10 
a = 8'd160; b = 8'd221;  #10 
a = 8'd160; b = 8'd222;  #10 
a = 8'd160; b = 8'd223;  #10 
a = 8'd160; b = 8'd224;  #10 
a = 8'd160; b = 8'd225;  #10 
a = 8'd160; b = 8'd226;  #10 
a = 8'd160; b = 8'd227;  #10 
a = 8'd160; b = 8'd228;  #10 
a = 8'd160; b = 8'd229;  #10 
a = 8'd160; b = 8'd230;  #10 
a = 8'd160; b = 8'd231;  #10 
a = 8'd160; b = 8'd232;  #10 
a = 8'd160; b = 8'd233;  #10 
a = 8'd160; b = 8'd234;  #10 
a = 8'd160; b = 8'd235;  #10 
a = 8'd160; b = 8'd236;  #10 
a = 8'd160; b = 8'd237;  #10 
a = 8'd160; b = 8'd238;  #10 
a = 8'd160; b = 8'd239;  #10 
a = 8'd160; b = 8'd240;  #10 
a = 8'd160; b = 8'd241;  #10 
a = 8'd160; b = 8'd242;  #10 
a = 8'd160; b = 8'd243;  #10 
a = 8'd160; b = 8'd244;  #10 
a = 8'd160; b = 8'd245;  #10 
a = 8'd160; b = 8'd246;  #10 
a = 8'd160; b = 8'd247;  #10 
a = 8'd160; b = 8'd248;  #10 
a = 8'd160; b = 8'd249;  #10 
a = 8'd160; b = 8'd250;  #10 
a = 8'd160; b = 8'd251;  #10 
a = 8'd160; b = 8'd252;  #10 
a = 8'd160; b = 8'd253;  #10 
a = 8'd160; b = 8'd254;  #10 
a = 8'd160; b = 8'd255;  #10 
a = 8'd161; b = 8'd0;  #10 
a = 8'd161; b = 8'd1;  #10 
a = 8'd161; b = 8'd2;  #10 
a = 8'd161; b = 8'd3;  #10 
a = 8'd161; b = 8'd4;  #10 
a = 8'd161; b = 8'd5;  #10 
a = 8'd161; b = 8'd6;  #10 
a = 8'd161; b = 8'd7;  #10 
a = 8'd161; b = 8'd8;  #10 
a = 8'd161; b = 8'd9;  #10 
a = 8'd161; b = 8'd10;  #10 
a = 8'd161; b = 8'd11;  #10 
a = 8'd161; b = 8'd12;  #10 
a = 8'd161; b = 8'd13;  #10 
a = 8'd161; b = 8'd14;  #10 
a = 8'd161; b = 8'd15;  #10 
a = 8'd161; b = 8'd16;  #10 
a = 8'd161; b = 8'd17;  #10 
a = 8'd161; b = 8'd18;  #10 
a = 8'd161; b = 8'd19;  #10 
a = 8'd161; b = 8'd20;  #10 
a = 8'd161; b = 8'd21;  #10 
a = 8'd161; b = 8'd22;  #10 
a = 8'd161; b = 8'd23;  #10 
a = 8'd161; b = 8'd24;  #10 
a = 8'd161; b = 8'd25;  #10 
a = 8'd161; b = 8'd26;  #10 
a = 8'd161; b = 8'd27;  #10 
a = 8'd161; b = 8'd28;  #10 
a = 8'd161; b = 8'd29;  #10 
a = 8'd161; b = 8'd30;  #10 
a = 8'd161; b = 8'd31;  #10 
a = 8'd161; b = 8'd32;  #10 
a = 8'd161; b = 8'd33;  #10 
a = 8'd161; b = 8'd34;  #10 
a = 8'd161; b = 8'd35;  #10 
a = 8'd161; b = 8'd36;  #10 
a = 8'd161; b = 8'd37;  #10 
a = 8'd161; b = 8'd38;  #10 
a = 8'd161; b = 8'd39;  #10 
a = 8'd161; b = 8'd40;  #10 
a = 8'd161; b = 8'd41;  #10 
a = 8'd161; b = 8'd42;  #10 
a = 8'd161; b = 8'd43;  #10 
a = 8'd161; b = 8'd44;  #10 
a = 8'd161; b = 8'd45;  #10 
a = 8'd161; b = 8'd46;  #10 
a = 8'd161; b = 8'd47;  #10 
a = 8'd161; b = 8'd48;  #10 
a = 8'd161; b = 8'd49;  #10 
a = 8'd161; b = 8'd50;  #10 
a = 8'd161; b = 8'd51;  #10 
a = 8'd161; b = 8'd52;  #10 
a = 8'd161; b = 8'd53;  #10 
a = 8'd161; b = 8'd54;  #10 
a = 8'd161; b = 8'd55;  #10 
a = 8'd161; b = 8'd56;  #10 
a = 8'd161; b = 8'd57;  #10 
a = 8'd161; b = 8'd58;  #10 
a = 8'd161; b = 8'd59;  #10 
a = 8'd161; b = 8'd60;  #10 
a = 8'd161; b = 8'd61;  #10 
a = 8'd161; b = 8'd62;  #10 
a = 8'd161; b = 8'd63;  #10 
a = 8'd161; b = 8'd64;  #10 
a = 8'd161; b = 8'd65;  #10 
a = 8'd161; b = 8'd66;  #10 
a = 8'd161; b = 8'd67;  #10 
a = 8'd161; b = 8'd68;  #10 
a = 8'd161; b = 8'd69;  #10 
a = 8'd161; b = 8'd70;  #10 
a = 8'd161; b = 8'd71;  #10 
a = 8'd161; b = 8'd72;  #10 
a = 8'd161; b = 8'd73;  #10 
a = 8'd161; b = 8'd74;  #10 
a = 8'd161; b = 8'd75;  #10 
a = 8'd161; b = 8'd76;  #10 
a = 8'd161; b = 8'd77;  #10 
a = 8'd161; b = 8'd78;  #10 
a = 8'd161; b = 8'd79;  #10 
a = 8'd161; b = 8'd80;  #10 
a = 8'd161; b = 8'd81;  #10 
a = 8'd161; b = 8'd82;  #10 
a = 8'd161; b = 8'd83;  #10 
a = 8'd161; b = 8'd84;  #10 
a = 8'd161; b = 8'd85;  #10 
a = 8'd161; b = 8'd86;  #10 
a = 8'd161; b = 8'd87;  #10 
a = 8'd161; b = 8'd88;  #10 
a = 8'd161; b = 8'd89;  #10 
a = 8'd161; b = 8'd90;  #10 
a = 8'd161; b = 8'd91;  #10 
a = 8'd161; b = 8'd92;  #10 
a = 8'd161; b = 8'd93;  #10 
a = 8'd161; b = 8'd94;  #10 
a = 8'd161; b = 8'd95;  #10 
a = 8'd161; b = 8'd96;  #10 
a = 8'd161; b = 8'd97;  #10 
a = 8'd161; b = 8'd98;  #10 
a = 8'd161; b = 8'd99;  #10 
a = 8'd161; b = 8'd100;  #10 
a = 8'd161; b = 8'd101;  #10 
a = 8'd161; b = 8'd102;  #10 
a = 8'd161; b = 8'd103;  #10 
a = 8'd161; b = 8'd104;  #10 
a = 8'd161; b = 8'd105;  #10 
a = 8'd161; b = 8'd106;  #10 
a = 8'd161; b = 8'd107;  #10 
a = 8'd161; b = 8'd108;  #10 
a = 8'd161; b = 8'd109;  #10 
a = 8'd161; b = 8'd110;  #10 
a = 8'd161; b = 8'd111;  #10 
a = 8'd161; b = 8'd112;  #10 
a = 8'd161; b = 8'd113;  #10 
a = 8'd161; b = 8'd114;  #10 
a = 8'd161; b = 8'd115;  #10 
a = 8'd161; b = 8'd116;  #10 
a = 8'd161; b = 8'd117;  #10 
a = 8'd161; b = 8'd118;  #10 
a = 8'd161; b = 8'd119;  #10 
a = 8'd161; b = 8'd120;  #10 
a = 8'd161; b = 8'd121;  #10 
a = 8'd161; b = 8'd122;  #10 
a = 8'd161; b = 8'd123;  #10 
a = 8'd161; b = 8'd124;  #10 
a = 8'd161; b = 8'd125;  #10 
a = 8'd161; b = 8'd126;  #10 
a = 8'd161; b = 8'd127;  #10 
a = 8'd161; b = 8'd128;  #10 
a = 8'd161; b = 8'd129;  #10 
a = 8'd161; b = 8'd130;  #10 
a = 8'd161; b = 8'd131;  #10 
a = 8'd161; b = 8'd132;  #10 
a = 8'd161; b = 8'd133;  #10 
a = 8'd161; b = 8'd134;  #10 
a = 8'd161; b = 8'd135;  #10 
a = 8'd161; b = 8'd136;  #10 
a = 8'd161; b = 8'd137;  #10 
a = 8'd161; b = 8'd138;  #10 
a = 8'd161; b = 8'd139;  #10 
a = 8'd161; b = 8'd140;  #10 
a = 8'd161; b = 8'd141;  #10 
a = 8'd161; b = 8'd142;  #10 
a = 8'd161; b = 8'd143;  #10 
a = 8'd161; b = 8'd144;  #10 
a = 8'd161; b = 8'd145;  #10 
a = 8'd161; b = 8'd146;  #10 
a = 8'd161; b = 8'd147;  #10 
a = 8'd161; b = 8'd148;  #10 
a = 8'd161; b = 8'd149;  #10 
a = 8'd161; b = 8'd150;  #10 
a = 8'd161; b = 8'd151;  #10 
a = 8'd161; b = 8'd152;  #10 
a = 8'd161; b = 8'd153;  #10 
a = 8'd161; b = 8'd154;  #10 
a = 8'd161; b = 8'd155;  #10 
a = 8'd161; b = 8'd156;  #10 
a = 8'd161; b = 8'd157;  #10 
a = 8'd161; b = 8'd158;  #10 
a = 8'd161; b = 8'd159;  #10 
a = 8'd161; b = 8'd160;  #10 
a = 8'd161; b = 8'd161;  #10 
a = 8'd161; b = 8'd162;  #10 
a = 8'd161; b = 8'd163;  #10 
a = 8'd161; b = 8'd164;  #10 
a = 8'd161; b = 8'd165;  #10 
a = 8'd161; b = 8'd166;  #10 
a = 8'd161; b = 8'd167;  #10 
a = 8'd161; b = 8'd168;  #10 
a = 8'd161; b = 8'd169;  #10 
a = 8'd161; b = 8'd170;  #10 
a = 8'd161; b = 8'd171;  #10 
a = 8'd161; b = 8'd172;  #10 
a = 8'd161; b = 8'd173;  #10 
a = 8'd161; b = 8'd174;  #10 
a = 8'd161; b = 8'd175;  #10 
a = 8'd161; b = 8'd176;  #10 
a = 8'd161; b = 8'd177;  #10 
a = 8'd161; b = 8'd178;  #10 
a = 8'd161; b = 8'd179;  #10 
a = 8'd161; b = 8'd180;  #10 
a = 8'd161; b = 8'd181;  #10 
a = 8'd161; b = 8'd182;  #10 
a = 8'd161; b = 8'd183;  #10 
a = 8'd161; b = 8'd184;  #10 
a = 8'd161; b = 8'd185;  #10 
a = 8'd161; b = 8'd186;  #10 
a = 8'd161; b = 8'd187;  #10 
a = 8'd161; b = 8'd188;  #10 
a = 8'd161; b = 8'd189;  #10 
a = 8'd161; b = 8'd190;  #10 
a = 8'd161; b = 8'd191;  #10 
a = 8'd161; b = 8'd192;  #10 
a = 8'd161; b = 8'd193;  #10 
a = 8'd161; b = 8'd194;  #10 
a = 8'd161; b = 8'd195;  #10 
a = 8'd161; b = 8'd196;  #10 
a = 8'd161; b = 8'd197;  #10 
a = 8'd161; b = 8'd198;  #10 
a = 8'd161; b = 8'd199;  #10 
a = 8'd161; b = 8'd200;  #10 
a = 8'd161; b = 8'd201;  #10 
a = 8'd161; b = 8'd202;  #10 
a = 8'd161; b = 8'd203;  #10 
a = 8'd161; b = 8'd204;  #10 
a = 8'd161; b = 8'd205;  #10 
a = 8'd161; b = 8'd206;  #10 
a = 8'd161; b = 8'd207;  #10 
a = 8'd161; b = 8'd208;  #10 
a = 8'd161; b = 8'd209;  #10 
a = 8'd161; b = 8'd210;  #10 
a = 8'd161; b = 8'd211;  #10 
a = 8'd161; b = 8'd212;  #10 
a = 8'd161; b = 8'd213;  #10 
a = 8'd161; b = 8'd214;  #10 
a = 8'd161; b = 8'd215;  #10 
a = 8'd161; b = 8'd216;  #10 
a = 8'd161; b = 8'd217;  #10 
a = 8'd161; b = 8'd218;  #10 
a = 8'd161; b = 8'd219;  #10 
a = 8'd161; b = 8'd220;  #10 
a = 8'd161; b = 8'd221;  #10 
a = 8'd161; b = 8'd222;  #10 
a = 8'd161; b = 8'd223;  #10 
a = 8'd161; b = 8'd224;  #10 
a = 8'd161; b = 8'd225;  #10 
a = 8'd161; b = 8'd226;  #10 
a = 8'd161; b = 8'd227;  #10 
a = 8'd161; b = 8'd228;  #10 
a = 8'd161; b = 8'd229;  #10 
a = 8'd161; b = 8'd230;  #10 
a = 8'd161; b = 8'd231;  #10 
a = 8'd161; b = 8'd232;  #10 
a = 8'd161; b = 8'd233;  #10 
a = 8'd161; b = 8'd234;  #10 
a = 8'd161; b = 8'd235;  #10 
a = 8'd161; b = 8'd236;  #10 
a = 8'd161; b = 8'd237;  #10 
a = 8'd161; b = 8'd238;  #10 
a = 8'd161; b = 8'd239;  #10 
a = 8'd161; b = 8'd240;  #10 
a = 8'd161; b = 8'd241;  #10 
a = 8'd161; b = 8'd242;  #10 
a = 8'd161; b = 8'd243;  #10 
a = 8'd161; b = 8'd244;  #10 
a = 8'd161; b = 8'd245;  #10 
a = 8'd161; b = 8'd246;  #10 
a = 8'd161; b = 8'd247;  #10 
a = 8'd161; b = 8'd248;  #10 
a = 8'd161; b = 8'd249;  #10 
a = 8'd161; b = 8'd250;  #10 
a = 8'd161; b = 8'd251;  #10 
a = 8'd161; b = 8'd252;  #10 
a = 8'd161; b = 8'd253;  #10 
a = 8'd161; b = 8'd254;  #10 
a = 8'd161; b = 8'd255;  #10 
a = 8'd162; b = 8'd0;  #10 
a = 8'd162; b = 8'd1;  #10 
a = 8'd162; b = 8'd2;  #10 
a = 8'd162; b = 8'd3;  #10 
a = 8'd162; b = 8'd4;  #10 
a = 8'd162; b = 8'd5;  #10 
a = 8'd162; b = 8'd6;  #10 
a = 8'd162; b = 8'd7;  #10 
a = 8'd162; b = 8'd8;  #10 
a = 8'd162; b = 8'd9;  #10 
a = 8'd162; b = 8'd10;  #10 
a = 8'd162; b = 8'd11;  #10 
a = 8'd162; b = 8'd12;  #10 
a = 8'd162; b = 8'd13;  #10 
a = 8'd162; b = 8'd14;  #10 
a = 8'd162; b = 8'd15;  #10 
a = 8'd162; b = 8'd16;  #10 
a = 8'd162; b = 8'd17;  #10 
a = 8'd162; b = 8'd18;  #10 
a = 8'd162; b = 8'd19;  #10 
a = 8'd162; b = 8'd20;  #10 
a = 8'd162; b = 8'd21;  #10 
a = 8'd162; b = 8'd22;  #10 
a = 8'd162; b = 8'd23;  #10 
a = 8'd162; b = 8'd24;  #10 
a = 8'd162; b = 8'd25;  #10 
a = 8'd162; b = 8'd26;  #10 
a = 8'd162; b = 8'd27;  #10 
a = 8'd162; b = 8'd28;  #10 
a = 8'd162; b = 8'd29;  #10 
a = 8'd162; b = 8'd30;  #10 
a = 8'd162; b = 8'd31;  #10 
a = 8'd162; b = 8'd32;  #10 
a = 8'd162; b = 8'd33;  #10 
a = 8'd162; b = 8'd34;  #10 
a = 8'd162; b = 8'd35;  #10 
a = 8'd162; b = 8'd36;  #10 
a = 8'd162; b = 8'd37;  #10 
a = 8'd162; b = 8'd38;  #10 
a = 8'd162; b = 8'd39;  #10 
a = 8'd162; b = 8'd40;  #10 
a = 8'd162; b = 8'd41;  #10 
a = 8'd162; b = 8'd42;  #10 
a = 8'd162; b = 8'd43;  #10 
a = 8'd162; b = 8'd44;  #10 
a = 8'd162; b = 8'd45;  #10 
a = 8'd162; b = 8'd46;  #10 
a = 8'd162; b = 8'd47;  #10 
a = 8'd162; b = 8'd48;  #10 
a = 8'd162; b = 8'd49;  #10 
a = 8'd162; b = 8'd50;  #10 
a = 8'd162; b = 8'd51;  #10 
a = 8'd162; b = 8'd52;  #10 
a = 8'd162; b = 8'd53;  #10 
a = 8'd162; b = 8'd54;  #10 
a = 8'd162; b = 8'd55;  #10 
a = 8'd162; b = 8'd56;  #10 
a = 8'd162; b = 8'd57;  #10 
a = 8'd162; b = 8'd58;  #10 
a = 8'd162; b = 8'd59;  #10 
a = 8'd162; b = 8'd60;  #10 
a = 8'd162; b = 8'd61;  #10 
a = 8'd162; b = 8'd62;  #10 
a = 8'd162; b = 8'd63;  #10 
a = 8'd162; b = 8'd64;  #10 
a = 8'd162; b = 8'd65;  #10 
a = 8'd162; b = 8'd66;  #10 
a = 8'd162; b = 8'd67;  #10 
a = 8'd162; b = 8'd68;  #10 
a = 8'd162; b = 8'd69;  #10 
a = 8'd162; b = 8'd70;  #10 
a = 8'd162; b = 8'd71;  #10 
a = 8'd162; b = 8'd72;  #10 
a = 8'd162; b = 8'd73;  #10 
a = 8'd162; b = 8'd74;  #10 
a = 8'd162; b = 8'd75;  #10 
a = 8'd162; b = 8'd76;  #10 
a = 8'd162; b = 8'd77;  #10 
a = 8'd162; b = 8'd78;  #10 
a = 8'd162; b = 8'd79;  #10 
a = 8'd162; b = 8'd80;  #10 
a = 8'd162; b = 8'd81;  #10 
a = 8'd162; b = 8'd82;  #10 
a = 8'd162; b = 8'd83;  #10 
a = 8'd162; b = 8'd84;  #10 
a = 8'd162; b = 8'd85;  #10 
a = 8'd162; b = 8'd86;  #10 
a = 8'd162; b = 8'd87;  #10 
a = 8'd162; b = 8'd88;  #10 
a = 8'd162; b = 8'd89;  #10 
a = 8'd162; b = 8'd90;  #10 
a = 8'd162; b = 8'd91;  #10 
a = 8'd162; b = 8'd92;  #10 
a = 8'd162; b = 8'd93;  #10 
a = 8'd162; b = 8'd94;  #10 
a = 8'd162; b = 8'd95;  #10 
a = 8'd162; b = 8'd96;  #10 
a = 8'd162; b = 8'd97;  #10 
a = 8'd162; b = 8'd98;  #10 
a = 8'd162; b = 8'd99;  #10 
a = 8'd162; b = 8'd100;  #10 
a = 8'd162; b = 8'd101;  #10 
a = 8'd162; b = 8'd102;  #10 
a = 8'd162; b = 8'd103;  #10 
a = 8'd162; b = 8'd104;  #10 
a = 8'd162; b = 8'd105;  #10 
a = 8'd162; b = 8'd106;  #10 
a = 8'd162; b = 8'd107;  #10 
a = 8'd162; b = 8'd108;  #10 
a = 8'd162; b = 8'd109;  #10 
a = 8'd162; b = 8'd110;  #10 
a = 8'd162; b = 8'd111;  #10 
a = 8'd162; b = 8'd112;  #10 
a = 8'd162; b = 8'd113;  #10 
a = 8'd162; b = 8'd114;  #10 
a = 8'd162; b = 8'd115;  #10 
a = 8'd162; b = 8'd116;  #10 
a = 8'd162; b = 8'd117;  #10 
a = 8'd162; b = 8'd118;  #10 
a = 8'd162; b = 8'd119;  #10 
a = 8'd162; b = 8'd120;  #10 
a = 8'd162; b = 8'd121;  #10 
a = 8'd162; b = 8'd122;  #10 
a = 8'd162; b = 8'd123;  #10 
a = 8'd162; b = 8'd124;  #10 
a = 8'd162; b = 8'd125;  #10 
a = 8'd162; b = 8'd126;  #10 
a = 8'd162; b = 8'd127;  #10 
a = 8'd162; b = 8'd128;  #10 
a = 8'd162; b = 8'd129;  #10 
a = 8'd162; b = 8'd130;  #10 
a = 8'd162; b = 8'd131;  #10 
a = 8'd162; b = 8'd132;  #10 
a = 8'd162; b = 8'd133;  #10 
a = 8'd162; b = 8'd134;  #10 
a = 8'd162; b = 8'd135;  #10 
a = 8'd162; b = 8'd136;  #10 
a = 8'd162; b = 8'd137;  #10 
a = 8'd162; b = 8'd138;  #10 
a = 8'd162; b = 8'd139;  #10 
a = 8'd162; b = 8'd140;  #10 
a = 8'd162; b = 8'd141;  #10 
a = 8'd162; b = 8'd142;  #10 
a = 8'd162; b = 8'd143;  #10 
a = 8'd162; b = 8'd144;  #10 
a = 8'd162; b = 8'd145;  #10 
a = 8'd162; b = 8'd146;  #10 
a = 8'd162; b = 8'd147;  #10 
a = 8'd162; b = 8'd148;  #10 
a = 8'd162; b = 8'd149;  #10 
a = 8'd162; b = 8'd150;  #10 
a = 8'd162; b = 8'd151;  #10 
a = 8'd162; b = 8'd152;  #10 
a = 8'd162; b = 8'd153;  #10 
a = 8'd162; b = 8'd154;  #10 
a = 8'd162; b = 8'd155;  #10 
a = 8'd162; b = 8'd156;  #10 
a = 8'd162; b = 8'd157;  #10 
a = 8'd162; b = 8'd158;  #10 
a = 8'd162; b = 8'd159;  #10 
a = 8'd162; b = 8'd160;  #10 
a = 8'd162; b = 8'd161;  #10 
a = 8'd162; b = 8'd162;  #10 
a = 8'd162; b = 8'd163;  #10 
a = 8'd162; b = 8'd164;  #10 
a = 8'd162; b = 8'd165;  #10 
a = 8'd162; b = 8'd166;  #10 
a = 8'd162; b = 8'd167;  #10 
a = 8'd162; b = 8'd168;  #10 
a = 8'd162; b = 8'd169;  #10 
a = 8'd162; b = 8'd170;  #10 
a = 8'd162; b = 8'd171;  #10 
a = 8'd162; b = 8'd172;  #10 
a = 8'd162; b = 8'd173;  #10 
a = 8'd162; b = 8'd174;  #10 
a = 8'd162; b = 8'd175;  #10 
a = 8'd162; b = 8'd176;  #10 
a = 8'd162; b = 8'd177;  #10 
a = 8'd162; b = 8'd178;  #10 
a = 8'd162; b = 8'd179;  #10 
a = 8'd162; b = 8'd180;  #10 
a = 8'd162; b = 8'd181;  #10 
a = 8'd162; b = 8'd182;  #10 
a = 8'd162; b = 8'd183;  #10 
a = 8'd162; b = 8'd184;  #10 
a = 8'd162; b = 8'd185;  #10 
a = 8'd162; b = 8'd186;  #10 
a = 8'd162; b = 8'd187;  #10 
a = 8'd162; b = 8'd188;  #10 
a = 8'd162; b = 8'd189;  #10 
a = 8'd162; b = 8'd190;  #10 
a = 8'd162; b = 8'd191;  #10 
a = 8'd162; b = 8'd192;  #10 
a = 8'd162; b = 8'd193;  #10 
a = 8'd162; b = 8'd194;  #10 
a = 8'd162; b = 8'd195;  #10 
a = 8'd162; b = 8'd196;  #10 
a = 8'd162; b = 8'd197;  #10 
a = 8'd162; b = 8'd198;  #10 
a = 8'd162; b = 8'd199;  #10 
a = 8'd162; b = 8'd200;  #10 
a = 8'd162; b = 8'd201;  #10 
a = 8'd162; b = 8'd202;  #10 
a = 8'd162; b = 8'd203;  #10 
a = 8'd162; b = 8'd204;  #10 
a = 8'd162; b = 8'd205;  #10 
a = 8'd162; b = 8'd206;  #10 
a = 8'd162; b = 8'd207;  #10 
a = 8'd162; b = 8'd208;  #10 
a = 8'd162; b = 8'd209;  #10 
a = 8'd162; b = 8'd210;  #10 
a = 8'd162; b = 8'd211;  #10 
a = 8'd162; b = 8'd212;  #10 
a = 8'd162; b = 8'd213;  #10 
a = 8'd162; b = 8'd214;  #10 
a = 8'd162; b = 8'd215;  #10 
a = 8'd162; b = 8'd216;  #10 
a = 8'd162; b = 8'd217;  #10 
a = 8'd162; b = 8'd218;  #10 
a = 8'd162; b = 8'd219;  #10 
a = 8'd162; b = 8'd220;  #10 
a = 8'd162; b = 8'd221;  #10 
a = 8'd162; b = 8'd222;  #10 
a = 8'd162; b = 8'd223;  #10 
a = 8'd162; b = 8'd224;  #10 
a = 8'd162; b = 8'd225;  #10 
a = 8'd162; b = 8'd226;  #10 
a = 8'd162; b = 8'd227;  #10 
a = 8'd162; b = 8'd228;  #10 
a = 8'd162; b = 8'd229;  #10 
a = 8'd162; b = 8'd230;  #10 
a = 8'd162; b = 8'd231;  #10 
a = 8'd162; b = 8'd232;  #10 
a = 8'd162; b = 8'd233;  #10 
a = 8'd162; b = 8'd234;  #10 
a = 8'd162; b = 8'd235;  #10 
a = 8'd162; b = 8'd236;  #10 
a = 8'd162; b = 8'd237;  #10 
a = 8'd162; b = 8'd238;  #10 
a = 8'd162; b = 8'd239;  #10 
a = 8'd162; b = 8'd240;  #10 
a = 8'd162; b = 8'd241;  #10 
a = 8'd162; b = 8'd242;  #10 
a = 8'd162; b = 8'd243;  #10 
a = 8'd162; b = 8'd244;  #10 
a = 8'd162; b = 8'd245;  #10 
a = 8'd162; b = 8'd246;  #10 
a = 8'd162; b = 8'd247;  #10 
a = 8'd162; b = 8'd248;  #10 
a = 8'd162; b = 8'd249;  #10 
a = 8'd162; b = 8'd250;  #10 
a = 8'd162; b = 8'd251;  #10 
a = 8'd162; b = 8'd252;  #10 
a = 8'd162; b = 8'd253;  #10 
a = 8'd162; b = 8'd254;  #10 
a = 8'd162; b = 8'd255;  #10 
a = 8'd163; b = 8'd0;  #10 
a = 8'd163; b = 8'd1;  #10 
a = 8'd163; b = 8'd2;  #10 
a = 8'd163; b = 8'd3;  #10 
a = 8'd163; b = 8'd4;  #10 
a = 8'd163; b = 8'd5;  #10 
a = 8'd163; b = 8'd6;  #10 
a = 8'd163; b = 8'd7;  #10 
a = 8'd163; b = 8'd8;  #10 
a = 8'd163; b = 8'd9;  #10 
a = 8'd163; b = 8'd10;  #10 
a = 8'd163; b = 8'd11;  #10 
a = 8'd163; b = 8'd12;  #10 
a = 8'd163; b = 8'd13;  #10 
a = 8'd163; b = 8'd14;  #10 
a = 8'd163; b = 8'd15;  #10 
a = 8'd163; b = 8'd16;  #10 
a = 8'd163; b = 8'd17;  #10 
a = 8'd163; b = 8'd18;  #10 
a = 8'd163; b = 8'd19;  #10 
a = 8'd163; b = 8'd20;  #10 
a = 8'd163; b = 8'd21;  #10 
a = 8'd163; b = 8'd22;  #10 
a = 8'd163; b = 8'd23;  #10 
a = 8'd163; b = 8'd24;  #10 
a = 8'd163; b = 8'd25;  #10 
a = 8'd163; b = 8'd26;  #10 
a = 8'd163; b = 8'd27;  #10 
a = 8'd163; b = 8'd28;  #10 
a = 8'd163; b = 8'd29;  #10 
a = 8'd163; b = 8'd30;  #10 
a = 8'd163; b = 8'd31;  #10 
a = 8'd163; b = 8'd32;  #10 
a = 8'd163; b = 8'd33;  #10 
a = 8'd163; b = 8'd34;  #10 
a = 8'd163; b = 8'd35;  #10 
a = 8'd163; b = 8'd36;  #10 
a = 8'd163; b = 8'd37;  #10 
a = 8'd163; b = 8'd38;  #10 
a = 8'd163; b = 8'd39;  #10 
a = 8'd163; b = 8'd40;  #10 
a = 8'd163; b = 8'd41;  #10 
a = 8'd163; b = 8'd42;  #10 
a = 8'd163; b = 8'd43;  #10 
a = 8'd163; b = 8'd44;  #10 
a = 8'd163; b = 8'd45;  #10 
a = 8'd163; b = 8'd46;  #10 
a = 8'd163; b = 8'd47;  #10 
a = 8'd163; b = 8'd48;  #10 
a = 8'd163; b = 8'd49;  #10 
a = 8'd163; b = 8'd50;  #10 
a = 8'd163; b = 8'd51;  #10 
a = 8'd163; b = 8'd52;  #10 
a = 8'd163; b = 8'd53;  #10 
a = 8'd163; b = 8'd54;  #10 
a = 8'd163; b = 8'd55;  #10 
a = 8'd163; b = 8'd56;  #10 
a = 8'd163; b = 8'd57;  #10 
a = 8'd163; b = 8'd58;  #10 
a = 8'd163; b = 8'd59;  #10 
a = 8'd163; b = 8'd60;  #10 
a = 8'd163; b = 8'd61;  #10 
a = 8'd163; b = 8'd62;  #10 
a = 8'd163; b = 8'd63;  #10 
a = 8'd163; b = 8'd64;  #10 
a = 8'd163; b = 8'd65;  #10 
a = 8'd163; b = 8'd66;  #10 
a = 8'd163; b = 8'd67;  #10 
a = 8'd163; b = 8'd68;  #10 
a = 8'd163; b = 8'd69;  #10 
a = 8'd163; b = 8'd70;  #10 
a = 8'd163; b = 8'd71;  #10 
a = 8'd163; b = 8'd72;  #10 
a = 8'd163; b = 8'd73;  #10 
a = 8'd163; b = 8'd74;  #10 
a = 8'd163; b = 8'd75;  #10 
a = 8'd163; b = 8'd76;  #10 
a = 8'd163; b = 8'd77;  #10 
a = 8'd163; b = 8'd78;  #10 
a = 8'd163; b = 8'd79;  #10 
a = 8'd163; b = 8'd80;  #10 
a = 8'd163; b = 8'd81;  #10 
a = 8'd163; b = 8'd82;  #10 
a = 8'd163; b = 8'd83;  #10 
a = 8'd163; b = 8'd84;  #10 
a = 8'd163; b = 8'd85;  #10 
a = 8'd163; b = 8'd86;  #10 
a = 8'd163; b = 8'd87;  #10 
a = 8'd163; b = 8'd88;  #10 
a = 8'd163; b = 8'd89;  #10 
a = 8'd163; b = 8'd90;  #10 
a = 8'd163; b = 8'd91;  #10 
a = 8'd163; b = 8'd92;  #10 
a = 8'd163; b = 8'd93;  #10 
a = 8'd163; b = 8'd94;  #10 
a = 8'd163; b = 8'd95;  #10 
a = 8'd163; b = 8'd96;  #10 
a = 8'd163; b = 8'd97;  #10 
a = 8'd163; b = 8'd98;  #10 
a = 8'd163; b = 8'd99;  #10 
a = 8'd163; b = 8'd100;  #10 
a = 8'd163; b = 8'd101;  #10 
a = 8'd163; b = 8'd102;  #10 
a = 8'd163; b = 8'd103;  #10 
a = 8'd163; b = 8'd104;  #10 
a = 8'd163; b = 8'd105;  #10 
a = 8'd163; b = 8'd106;  #10 
a = 8'd163; b = 8'd107;  #10 
a = 8'd163; b = 8'd108;  #10 
a = 8'd163; b = 8'd109;  #10 
a = 8'd163; b = 8'd110;  #10 
a = 8'd163; b = 8'd111;  #10 
a = 8'd163; b = 8'd112;  #10 
a = 8'd163; b = 8'd113;  #10 
a = 8'd163; b = 8'd114;  #10 
a = 8'd163; b = 8'd115;  #10 
a = 8'd163; b = 8'd116;  #10 
a = 8'd163; b = 8'd117;  #10 
a = 8'd163; b = 8'd118;  #10 
a = 8'd163; b = 8'd119;  #10 
a = 8'd163; b = 8'd120;  #10 
a = 8'd163; b = 8'd121;  #10 
a = 8'd163; b = 8'd122;  #10 
a = 8'd163; b = 8'd123;  #10 
a = 8'd163; b = 8'd124;  #10 
a = 8'd163; b = 8'd125;  #10 
a = 8'd163; b = 8'd126;  #10 
a = 8'd163; b = 8'd127;  #10 
a = 8'd163; b = 8'd128;  #10 
a = 8'd163; b = 8'd129;  #10 
a = 8'd163; b = 8'd130;  #10 
a = 8'd163; b = 8'd131;  #10 
a = 8'd163; b = 8'd132;  #10 
a = 8'd163; b = 8'd133;  #10 
a = 8'd163; b = 8'd134;  #10 
a = 8'd163; b = 8'd135;  #10 
a = 8'd163; b = 8'd136;  #10 
a = 8'd163; b = 8'd137;  #10 
a = 8'd163; b = 8'd138;  #10 
a = 8'd163; b = 8'd139;  #10 
a = 8'd163; b = 8'd140;  #10 
a = 8'd163; b = 8'd141;  #10 
a = 8'd163; b = 8'd142;  #10 
a = 8'd163; b = 8'd143;  #10 
a = 8'd163; b = 8'd144;  #10 
a = 8'd163; b = 8'd145;  #10 
a = 8'd163; b = 8'd146;  #10 
a = 8'd163; b = 8'd147;  #10 
a = 8'd163; b = 8'd148;  #10 
a = 8'd163; b = 8'd149;  #10 
a = 8'd163; b = 8'd150;  #10 
a = 8'd163; b = 8'd151;  #10 
a = 8'd163; b = 8'd152;  #10 
a = 8'd163; b = 8'd153;  #10 
a = 8'd163; b = 8'd154;  #10 
a = 8'd163; b = 8'd155;  #10 
a = 8'd163; b = 8'd156;  #10 
a = 8'd163; b = 8'd157;  #10 
a = 8'd163; b = 8'd158;  #10 
a = 8'd163; b = 8'd159;  #10 
a = 8'd163; b = 8'd160;  #10 
a = 8'd163; b = 8'd161;  #10 
a = 8'd163; b = 8'd162;  #10 
a = 8'd163; b = 8'd163;  #10 
a = 8'd163; b = 8'd164;  #10 
a = 8'd163; b = 8'd165;  #10 
a = 8'd163; b = 8'd166;  #10 
a = 8'd163; b = 8'd167;  #10 
a = 8'd163; b = 8'd168;  #10 
a = 8'd163; b = 8'd169;  #10 
a = 8'd163; b = 8'd170;  #10 
a = 8'd163; b = 8'd171;  #10 
a = 8'd163; b = 8'd172;  #10 
a = 8'd163; b = 8'd173;  #10 
a = 8'd163; b = 8'd174;  #10 
a = 8'd163; b = 8'd175;  #10 
a = 8'd163; b = 8'd176;  #10 
a = 8'd163; b = 8'd177;  #10 
a = 8'd163; b = 8'd178;  #10 
a = 8'd163; b = 8'd179;  #10 
a = 8'd163; b = 8'd180;  #10 
a = 8'd163; b = 8'd181;  #10 
a = 8'd163; b = 8'd182;  #10 
a = 8'd163; b = 8'd183;  #10 
a = 8'd163; b = 8'd184;  #10 
a = 8'd163; b = 8'd185;  #10 
a = 8'd163; b = 8'd186;  #10 
a = 8'd163; b = 8'd187;  #10 
a = 8'd163; b = 8'd188;  #10 
a = 8'd163; b = 8'd189;  #10 
a = 8'd163; b = 8'd190;  #10 
a = 8'd163; b = 8'd191;  #10 
a = 8'd163; b = 8'd192;  #10 
a = 8'd163; b = 8'd193;  #10 
a = 8'd163; b = 8'd194;  #10 
a = 8'd163; b = 8'd195;  #10 
a = 8'd163; b = 8'd196;  #10 
a = 8'd163; b = 8'd197;  #10 
a = 8'd163; b = 8'd198;  #10 
a = 8'd163; b = 8'd199;  #10 
a = 8'd163; b = 8'd200;  #10 
a = 8'd163; b = 8'd201;  #10 
a = 8'd163; b = 8'd202;  #10 
a = 8'd163; b = 8'd203;  #10 
a = 8'd163; b = 8'd204;  #10 
a = 8'd163; b = 8'd205;  #10 
a = 8'd163; b = 8'd206;  #10 
a = 8'd163; b = 8'd207;  #10 
a = 8'd163; b = 8'd208;  #10 
a = 8'd163; b = 8'd209;  #10 
a = 8'd163; b = 8'd210;  #10 
a = 8'd163; b = 8'd211;  #10 
a = 8'd163; b = 8'd212;  #10 
a = 8'd163; b = 8'd213;  #10 
a = 8'd163; b = 8'd214;  #10 
a = 8'd163; b = 8'd215;  #10 
a = 8'd163; b = 8'd216;  #10 
a = 8'd163; b = 8'd217;  #10 
a = 8'd163; b = 8'd218;  #10 
a = 8'd163; b = 8'd219;  #10 
a = 8'd163; b = 8'd220;  #10 
a = 8'd163; b = 8'd221;  #10 
a = 8'd163; b = 8'd222;  #10 
a = 8'd163; b = 8'd223;  #10 
a = 8'd163; b = 8'd224;  #10 
a = 8'd163; b = 8'd225;  #10 
a = 8'd163; b = 8'd226;  #10 
a = 8'd163; b = 8'd227;  #10 
a = 8'd163; b = 8'd228;  #10 
a = 8'd163; b = 8'd229;  #10 
a = 8'd163; b = 8'd230;  #10 
a = 8'd163; b = 8'd231;  #10 
a = 8'd163; b = 8'd232;  #10 
a = 8'd163; b = 8'd233;  #10 
a = 8'd163; b = 8'd234;  #10 
a = 8'd163; b = 8'd235;  #10 
a = 8'd163; b = 8'd236;  #10 
a = 8'd163; b = 8'd237;  #10 
a = 8'd163; b = 8'd238;  #10 
a = 8'd163; b = 8'd239;  #10 
a = 8'd163; b = 8'd240;  #10 
a = 8'd163; b = 8'd241;  #10 
a = 8'd163; b = 8'd242;  #10 
a = 8'd163; b = 8'd243;  #10 
a = 8'd163; b = 8'd244;  #10 
a = 8'd163; b = 8'd245;  #10 
a = 8'd163; b = 8'd246;  #10 
a = 8'd163; b = 8'd247;  #10 
a = 8'd163; b = 8'd248;  #10 
a = 8'd163; b = 8'd249;  #10 
a = 8'd163; b = 8'd250;  #10 
a = 8'd163; b = 8'd251;  #10 
a = 8'd163; b = 8'd252;  #10 
a = 8'd163; b = 8'd253;  #10 
a = 8'd163; b = 8'd254;  #10 
a = 8'd163; b = 8'd255;  #10 
a = 8'd164; b = 8'd0;  #10 
a = 8'd164; b = 8'd1;  #10 
a = 8'd164; b = 8'd2;  #10 
a = 8'd164; b = 8'd3;  #10 
a = 8'd164; b = 8'd4;  #10 
a = 8'd164; b = 8'd5;  #10 
a = 8'd164; b = 8'd6;  #10 
a = 8'd164; b = 8'd7;  #10 
a = 8'd164; b = 8'd8;  #10 
a = 8'd164; b = 8'd9;  #10 
a = 8'd164; b = 8'd10;  #10 
a = 8'd164; b = 8'd11;  #10 
a = 8'd164; b = 8'd12;  #10 
a = 8'd164; b = 8'd13;  #10 
a = 8'd164; b = 8'd14;  #10 
a = 8'd164; b = 8'd15;  #10 
a = 8'd164; b = 8'd16;  #10 
a = 8'd164; b = 8'd17;  #10 
a = 8'd164; b = 8'd18;  #10 
a = 8'd164; b = 8'd19;  #10 
a = 8'd164; b = 8'd20;  #10 
a = 8'd164; b = 8'd21;  #10 
a = 8'd164; b = 8'd22;  #10 
a = 8'd164; b = 8'd23;  #10 
a = 8'd164; b = 8'd24;  #10 
a = 8'd164; b = 8'd25;  #10 
a = 8'd164; b = 8'd26;  #10 
a = 8'd164; b = 8'd27;  #10 
a = 8'd164; b = 8'd28;  #10 
a = 8'd164; b = 8'd29;  #10 
a = 8'd164; b = 8'd30;  #10 
a = 8'd164; b = 8'd31;  #10 
a = 8'd164; b = 8'd32;  #10 
a = 8'd164; b = 8'd33;  #10 
a = 8'd164; b = 8'd34;  #10 
a = 8'd164; b = 8'd35;  #10 
a = 8'd164; b = 8'd36;  #10 
a = 8'd164; b = 8'd37;  #10 
a = 8'd164; b = 8'd38;  #10 
a = 8'd164; b = 8'd39;  #10 
a = 8'd164; b = 8'd40;  #10 
a = 8'd164; b = 8'd41;  #10 
a = 8'd164; b = 8'd42;  #10 
a = 8'd164; b = 8'd43;  #10 
a = 8'd164; b = 8'd44;  #10 
a = 8'd164; b = 8'd45;  #10 
a = 8'd164; b = 8'd46;  #10 
a = 8'd164; b = 8'd47;  #10 
a = 8'd164; b = 8'd48;  #10 
a = 8'd164; b = 8'd49;  #10 
a = 8'd164; b = 8'd50;  #10 
a = 8'd164; b = 8'd51;  #10 
a = 8'd164; b = 8'd52;  #10 
a = 8'd164; b = 8'd53;  #10 
a = 8'd164; b = 8'd54;  #10 
a = 8'd164; b = 8'd55;  #10 
a = 8'd164; b = 8'd56;  #10 
a = 8'd164; b = 8'd57;  #10 
a = 8'd164; b = 8'd58;  #10 
a = 8'd164; b = 8'd59;  #10 
a = 8'd164; b = 8'd60;  #10 
a = 8'd164; b = 8'd61;  #10 
a = 8'd164; b = 8'd62;  #10 
a = 8'd164; b = 8'd63;  #10 
a = 8'd164; b = 8'd64;  #10 
a = 8'd164; b = 8'd65;  #10 
a = 8'd164; b = 8'd66;  #10 
a = 8'd164; b = 8'd67;  #10 
a = 8'd164; b = 8'd68;  #10 
a = 8'd164; b = 8'd69;  #10 
a = 8'd164; b = 8'd70;  #10 
a = 8'd164; b = 8'd71;  #10 
a = 8'd164; b = 8'd72;  #10 
a = 8'd164; b = 8'd73;  #10 
a = 8'd164; b = 8'd74;  #10 
a = 8'd164; b = 8'd75;  #10 
a = 8'd164; b = 8'd76;  #10 
a = 8'd164; b = 8'd77;  #10 
a = 8'd164; b = 8'd78;  #10 
a = 8'd164; b = 8'd79;  #10 
a = 8'd164; b = 8'd80;  #10 
a = 8'd164; b = 8'd81;  #10 
a = 8'd164; b = 8'd82;  #10 
a = 8'd164; b = 8'd83;  #10 
a = 8'd164; b = 8'd84;  #10 
a = 8'd164; b = 8'd85;  #10 
a = 8'd164; b = 8'd86;  #10 
a = 8'd164; b = 8'd87;  #10 
a = 8'd164; b = 8'd88;  #10 
a = 8'd164; b = 8'd89;  #10 
a = 8'd164; b = 8'd90;  #10 
a = 8'd164; b = 8'd91;  #10 
a = 8'd164; b = 8'd92;  #10 
a = 8'd164; b = 8'd93;  #10 
a = 8'd164; b = 8'd94;  #10 
a = 8'd164; b = 8'd95;  #10 
a = 8'd164; b = 8'd96;  #10 
a = 8'd164; b = 8'd97;  #10 
a = 8'd164; b = 8'd98;  #10 
a = 8'd164; b = 8'd99;  #10 
a = 8'd164; b = 8'd100;  #10 
a = 8'd164; b = 8'd101;  #10 
a = 8'd164; b = 8'd102;  #10 
a = 8'd164; b = 8'd103;  #10 
a = 8'd164; b = 8'd104;  #10 
a = 8'd164; b = 8'd105;  #10 
a = 8'd164; b = 8'd106;  #10 
a = 8'd164; b = 8'd107;  #10 
a = 8'd164; b = 8'd108;  #10 
a = 8'd164; b = 8'd109;  #10 
a = 8'd164; b = 8'd110;  #10 
a = 8'd164; b = 8'd111;  #10 
a = 8'd164; b = 8'd112;  #10 
a = 8'd164; b = 8'd113;  #10 
a = 8'd164; b = 8'd114;  #10 
a = 8'd164; b = 8'd115;  #10 
a = 8'd164; b = 8'd116;  #10 
a = 8'd164; b = 8'd117;  #10 
a = 8'd164; b = 8'd118;  #10 
a = 8'd164; b = 8'd119;  #10 
a = 8'd164; b = 8'd120;  #10 
a = 8'd164; b = 8'd121;  #10 
a = 8'd164; b = 8'd122;  #10 
a = 8'd164; b = 8'd123;  #10 
a = 8'd164; b = 8'd124;  #10 
a = 8'd164; b = 8'd125;  #10 
a = 8'd164; b = 8'd126;  #10 
a = 8'd164; b = 8'd127;  #10 
a = 8'd164; b = 8'd128;  #10 
a = 8'd164; b = 8'd129;  #10 
a = 8'd164; b = 8'd130;  #10 
a = 8'd164; b = 8'd131;  #10 
a = 8'd164; b = 8'd132;  #10 
a = 8'd164; b = 8'd133;  #10 
a = 8'd164; b = 8'd134;  #10 
a = 8'd164; b = 8'd135;  #10 
a = 8'd164; b = 8'd136;  #10 
a = 8'd164; b = 8'd137;  #10 
a = 8'd164; b = 8'd138;  #10 
a = 8'd164; b = 8'd139;  #10 
a = 8'd164; b = 8'd140;  #10 
a = 8'd164; b = 8'd141;  #10 
a = 8'd164; b = 8'd142;  #10 
a = 8'd164; b = 8'd143;  #10 
a = 8'd164; b = 8'd144;  #10 
a = 8'd164; b = 8'd145;  #10 
a = 8'd164; b = 8'd146;  #10 
a = 8'd164; b = 8'd147;  #10 
a = 8'd164; b = 8'd148;  #10 
a = 8'd164; b = 8'd149;  #10 
a = 8'd164; b = 8'd150;  #10 
a = 8'd164; b = 8'd151;  #10 
a = 8'd164; b = 8'd152;  #10 
a = 8'd164; b = 8'd153;  #10 
a = 8'd164; b = 8'd154;  #10 
a = 8'd164; b = 8'd155;  #10 
a = 8'd164; b = 8'd156;  #10 
a = 8'd164; b = 8'd157;  #10 
a = 8'd164; b = 8'd158;  #10 
a = 8'd164; b = 8'd159;  #10 
a = 8'd164; b = 8'd160;  #10 
a = 8'd164; b = 8'd161;  #10 
a = 8'd164; b = 8'd162;  #10 
a = 8'd164; b = 8'd163;  #10 
a = 8'd164; b = 8'd164;  #10 
a = 8'd164; b = 8'd165;  #10 
a = 8'd164; b = 8'd166;  #10 
a = 8'd164; b = 8'd167;  #10 
a = 8'd164; b = 8'd168;  #10 
a = 8'd164; b = 8'd169;  #10 
a = 8'd164; b = 8'd170;  #10 
a = 8'd164; b = 8'd171;  #10 
a = 8'd164; b = 8'd172;  #10 
a = 8'd164; b = 8'd173;  #10 
a = 8'd164; b = 8'd174;  #10 
a = 8'd164; b = 8'd175;  #10 
a = 8'd164; b = 8'd176;  #10 
a = 8'd164; b = 8'd177;  #10 
a = 8'd164; b = 8'd178;  #10 
a = 8'd164; b = 8'd179;  #10 
a = 8'd164; b = 8'd180;  #10 
a = 8'd164; b = 8'd181;  #10 
a = 8'd164; b = 8'd182;  #10 
a = 8'd164; b = 8'd183;  #10 
a = 8'd164; b = 8'd184;  #10 
a = 8'd164; b = 8'd185;  #10 
a = 8'd164; b = 8'd186;  #10 
a = 8'd164; b = 8'd187;  #10 
a = 8'd164; b = 8'd188;  #10 
a = 8'd164; b = 8'd189;  #10 
a = 8'd164; b = 8'd190;  #10 
a = 8'd164; b = 8'd191;  #10 
a = 8'd164; b = 8'd192;  #10 
a = 8'd164; b = 8'd193;  #10 
a = 8'd164; b = 8'd194;  #10 
a = 8'd164; b = 8'd195;  #10 
a = 8'd164; b = 8'd196;  #10 
a = 8'd164; b = 8'd197;  #10 
a = 8'd164; b = 8'd198;  #10 
a = 8'd164; b = 8'd199;  #10 
a = 8'd164; b = 8'd200;  #10 
a = 8'd164; b = 8'd201;  #10 
a = 8'd164; b = 8'd202;  #10 
a = 8'd164; b = 8'd203;  #10 
a = 8'd164; b = 8'd204;  #10 
a = 8'd164; b = 8'd205;  #10 
a = 8'd164; b = 8'd206;  #10 
a = 8'd164; b = 8'd207;  #10 
a = 8'd164; b = 8'd208;  #10 
a = 8'd164; b = 8'd209;  #10 
a = 8'd164; b = 8'd210;  #10 
a = 8'd164; b = 8'd211;  #10 
a = 8'd164; b = 8'd212;  #10 
a = 8'd164; b = 8'd213;  #10 
a = 8'd164; b = 8'd214;  #10 
a = 8'd164; b = 8'd215;  #10 
a = 8'd164; b = 8'd216;  #10 
a = 8'd164; b = 8'd217;  #10 
a = 8'd164; b = 8'd218;  #10 
a = 8'd164; b = 8'd219;  #10 
a = 8'd164; b = 8'd220;  #10 
a = 8'd164; b = 8'd221;  #10 
a = 8'd164; b = 8'd222;  #10 
a = 8'd164; b = 8'd223;  #10 
a = 8'd164; b = 8'd224;  #10 
a = 8'd164; b = 8'd225;  #10 
a = 8'd164; b = 8'd226;  #10 
a = 8'd164; b = 8'd227;  #10 
a = 8'd164; b = 8'd228;  #10 
a = 8'd164; b = 8'd229;  #10 
a = 8'd164; b = 8'd230;  #10 
a = 8'd164; b = 8'd231;  #10 
a = 8'd164; b = 8'd232;  #10 
a = 8'd164; b = 8'd233;  #10 
a = 8'd164; b = 8'd234;  #10 
a = 8'd164; b = 8'd235;  #10 
a = 8'd164; b = 8'd236;  #10 
a = 8'd164; b = 8'd237;  #10 
a = 8'd164; b = 8'd238;  #10 
a = 8'd164; b = 8'd239;  #10 
a = 8'd164; b = 8'd240;  #10 
a = 8'd164; b = 8'd241;  #10 
a = 8'd164; b = 8'd242;  #10 
a = 8'd164; b = 8'd243;  #10 
a = 8'd164; b = 8'd244;  #10 
a = 8'd164; b = 8'd245;  #10 
a = 8'd164; b = 8'd246;  #10 
a = 8'd164; b = 8'd247;  #10 
a = 8'd164; b = 8'd248;  #10 
a = 8'd164; b = 8'd249;  #10 
a = 8'd164; b = 8'd250;  #10 
a = 8'd164; b = 8'd251;  #10 
a = 8'd164; b = 8'd252;  #10 
a = 8'd164; b = 8'd253;  #10 
a = 8'd164; b = 8'd254;  #10 
a = 8'd164; b = 8'd255;  #10 
a = 8'd165; b = 8'd0;  #10 
a = 8'd165; b = 8'd1;  #10 
a = 8'd165; b = 8'd2;  #10 
a = 8'd165; b = 8'd3;  #10 
a = 8'd165; b = 8'd4;  #10 
a = 8'd165; b = 8'd5;  #10 
a = 8'd165; b = 8'd6;  #10 
a = 8'd165; b = 8'd7;  #10 
a = 8'd165; b = 8'd8;  #10 
a = 8'd165; b = 8'd9;  #10 
a = 8'd165; b = 8'd10;  #10 
a = 8'd165; b = 8'd11;  #10 
a = 8'd165; b = 8'd12;  #10 
a = 8'd165; b = 8'd13;  #10 
a = 8'd165; b = 8'd14;  #10 
a = 8'd165; b = 8'd15;  #10 
a = 8'd165; b = 8'd16;  #10 
a = 8'd165; b = 8'd17;  #10 
a = 8'd165; b = 8'd18;  #10 
a = 8'd165; b = 8'd19;  #10 
a = 8'd165; b = 8'd20;  #10 
a = 8'd165; b = 8'd21;  #10 
a = 8'd165; b = 8'd22;  #10 
a = 8'd165; b = 8'd23;  #10 
a = 8'd165; b = 8'd24;  #10 
a = 8'd165; b = 8'd25;  #10 
a = 8'd165; b = 8'd26;  #10 
a = 8'd165; b = 8'd27;  #10 
a = 8'd165; b = 8'd28;  #10 
a = 8'd165; b = 8'd29;  #10 
a = 8'd165; b = 8'd30;  #10 
a = 8'd165; b = 8'd31;  #10 
a = 8'd165; b = 8'd32;  #10 
a = 8'd165; b = 8'd33;  #10 
a = 8'd165; b = 8'd34;  #10 
a = 8'd165; b = 8'd35;  #10 
a = 8'd165; b = 8'd36;  #10 
a = 8'd165; b = 8'd37;  #10 
a = 8'd165; b = 8'd38;  #10 
a = 8'd165; b = 8'd39;  #10 
a = 8'd165; b = 8'd40;  #10 
a = 8'd165; b = 8'd41;  #10 
a = 8'd165; b = 8'd42;  #10 
a = 8'd165; b = 8'd43;  #10 
a = 8'd165; b = 8'd44;  #10 
a = 8'd165; b = 8'd45;  #10 
a = 8'd165; b = 8'd46;  #10 
a = 8'd165; b = 8'd47;  #10 
a = 8'd165; b = 8'd48;  #10 
a = 8'd165; b = 8'd49;  #10 
a = 8'd165; b = 8'd50;  #10 
a = 8'd165; b = 8'd51;  #10 
a = 8'd165; b = 8'd52;  #10 
a = 8'd165; b = 8'd53;  #10 
a = 8'd165; b = 8'd54;  #10 
a = 8'd165; b = 8'd55;  #10 
a = 8'd165; b = 8'd56;  #10 
a = 8'd165; b = 8'd57;  #10 
a = 8'd165; b = 8'd58;  #10 
a = 8'd165; b = 8'd59;  #10 
a = 8'd165; b = 8'd60;  #10 
a = 8'd165; b = 8'd61;  #10 
a = 8'd165; b = 8'd62;  #10 
a = 8'd165; b = 8'd63;  #10 
a = 8'd165; b = 8'd64;  #10 
a = 8'd165; b = 8'd65;  #10 
a = 8'd165; b = 8'd66;  #10 
a = 8'd165; b = 8'd67;  #10 
a = 8'd165; b = 8'd68;  #10 
a = 8'd165; b = 8'd69;  #10 
a = 8'd165; b = 8'd70;  #10 
a = 8'd165; b = 8'd71;  #10 
a = 8'd165; b = 8'd72;  #10 
a = 8'd165; b = 8'd73;  #10 
a = 8'd165; b = 8'd74;  #10 
a = 8'd165; b = 8'd75;  #10 
a = 8'd165; b = 8'd76;  #10 
a = 8'd165; b = 8'd77;  #10 
a = 8'd165; b = 8'd78;  #10 
a = 8'd165; b = 8'd79;  #10 
a = 8'd165; b = 8'd80;  #10 
a = 8'd165; b = 8'd81;  #10 
a = 8'd165; b = 8'd82;  #10 
a = 8'd165; b = 8'd83;  #10 
a = 8'd165; b = 8'd84;  #10 
a = 8'd165; b = 8'd85;  #10 
a = 8'd165; b = 8'd86;  #10 
a = 8'd165; b = 8'd87;  #10 
a = 8'd165; b = 8'd88;  #10 
a = 8'd165; b = 8'd89;  #10 
a = 8'd165; b = 8'd90;  #10 
a = 8'd165; b = 8'd91;  #10 
a = 8'd165; b = 8'd92;  #10 
a = 8'd165; b = 8'd93;  #10 
a = 8'd165; b = 8'd94;  #10 
a = 8'd165; b = 8'd95;  #10 
a = 8'd165; b = 8'd96;  #10 
a = 8'd165; b = 8'd97;  #10 
a = 8'd165; b = 8'd98;  #10 
a = 8'd165; b = 8'd99;  #10 
a = 8'd165; b = 8'd100;  #10 
a = 8'd165; b = 8'd101;  #10 
a = 8'd165; b = 8'd102;  #10 
a = 8'd165; b = 8'd103;  #10 
a = 8'd165; b = 8'd104;  #10 
a = 8'd165; b = 8'd105;  #10 
a = 8'd165; b = 8'd106;  #10 
a = 8'd165; b = 8'd107;  #10 
a = 8'd165; b = 8'd108;  #10 
a = 8'd165; b = 8'd109;  #10 
a = 8'd165; b = 8'd110;  #10 
a = 8'd165; b = 8'd111;  #10 
a = 8'd165; b = 8'd112;  #10 
a = 8'd165; b = 8'd113;  #10 
a = 8'd165; b = 8'd114;  #10 
a = 8'd165; b = 8'd115;  #10 
a = 8'd165; b = 8'd116;  #10 
a = 8'd165; b = 8'd117;  #10 
a = 8'd165; b = 8'd118;  #10 
a = 8'd165; b = 8'd119;  #10 
a = 8'd165; b = 8'd120;  #10 
a = 8'd165; b = 8'd121;  #10 
a = 8'd165; b = 8'd122;  #10 
a = 8'd165; b = 8'd123;  #10 
a = 8'd165; b = 8'd124;  #10 
a = 8'd165; b = 8'd125;  #10 
a = 8'd165; b = 8'd126;  #10 
a = 8'd165; b = 8'd127;  #10 
a = 8'd165; b = 8'd128;  #10 
a = 8'd165; b = 8'd129;  #10 
a = 8'd165; b = 8'd130;  #10 
a = 8'd165; b = 8'd131;  #10 
a = 8'd165; b = 8'd132;  #10 
a = 8'd165; b = 8'd133;  #10 
a = 8'd165; b = 8'd134;  #10 
a = 8'd165; b = 8'd135;  #10 
a = 8'd165; b = 8'd136;  #10 
a = 8'd165; b = 8'd137;  #10 
a = 8'd165; b = 8'd138;  #10 
a = 8'd165; b = 8'd139;  #10 
a = 8'd165; b = 8'd140;  #10 
a = 8'd165; b = 8'd141;  #10 
a = 8'd165; b = 8'd142;  #10 
a = 8'd165; b = 8'd143;  #10 
a = 8'd165; b = 8'd144;  #10 
a = 8'd165; b = 8'd145;  #10 
a = 8'd165; b = 8'd146;  #10 
a = 8'd165; b = 8'd147;  #10 
a = 8'd165; b = 8'd148;  #10 
a = 8'd165; b = 8'd149;  #10 
a = 8'd165; b = 8'd150;  #10 
a = 8'd165; b = 8'd151;  #10 
a = 8'd165; b = 8'd152;  #10 
a = 8'd165; b = 8'd153;  #10 
a = 8'd165; b = 8'd154;  #10 
a = 8'd165; b = 8'd155;  #10 
a = 8'd165; b = 8'd156;  #10 
a = 8'd165; b = 8'd157;  #10 
a = 8'd165; b = 8'd158;  #10 
a = 8'd165; b = 8'd159;  #10 
a = 8'd165; b = 8'd160;  #10 
a = 8'd165; b = 8'd161;  #10 
a = 8'd165; b = 8'd162;  #10 
a = 8'd165; b = 8'd163;  #10 
a = 8'd165; b = 8'd164;  #10 
a = 8'd165; b = 8'd165;  #10 
a = 8'd165; b = 8'd166;  #10 
a = 8'd165; b = 8'd167;  #10 
a = 8'd165; b = 8'd168;  #10 
a = 8'd165; b = 8'd169;  #10 
a = 8'd165; b = 8'd170;  #10 
a = 8'd165; b = 8'd171;  #10 
a = 8'd165; b = 8'd172;  #10 
a = 8'd165; b = 8'd173;  #10 
a = 8'd165; b = 8'd174;  #10 
a = 8'd165; b = 8'd175;  #10 
a = 8'd165; b = 8'd176;  #10 
a = 8'd165; b = 8'd177;  #10 
a = 8'd165; b = 8'd178;  #10 
a = 8'd165; b = 8'd179;  #10 
a = 8'd165; b = 8'd180;  #10 
a = 8'd165; b = 8'd181;  #10 
a = 8'd165; b = 8'd182;  #10 
a = 8'd165; b = 8'd183;  #10 
a = 8'd165; b = 8'd184;  #10 
a = 8'd165; b = 8'd185;  #10 
a = 8'd165; b = 8'd186;  #10 
a = 8'd165; b = 8'd187;  #10 
a = 8'd165; b = 8'd188;  #10 
a = 8'd165; b = 8'd189;  #10 
a = 8'd165; b = 8'd190;  #10 
a = 8'd165; b = 8'd191;  #10 
a = 8'd165; b = 8'd192;  #10 
a = 8'd165; b = 8'd193;  #10 
a = 8'd165; b = 8'd194;  #10 
a = 8'd165; b = 8'd195;  #10 
a = 8'd165; b = 8'd196;  #10 
a = 8'd165; b = 8'd197;  #10 
a = 8'd165; b = 8'd198;  #10 
a = 8'd165; b = 8'd199;  #10 
a = 8'd165; b = 8'd200;  #10 
a = 8'd165; b = 8'd201;  #10 
a = 8'd165; b = 8'd202;  #10 
a = 8'd165; b = 8'd203;  #10 
a = 8'd165; b = 8'd204;  #10 
a = 8'd165; b = 8'd205;  #10 
a = 8'd165; b = 8'd206;  #10 
a = 8'd165; b = 8'd207;  #10 
a = 8'd165; b = 8'd208;  #10 
a = 8'd165; b = 8'd209;  #10 
a = 8'd165; b = 8'd210;  #10 
a = 8'd165; b = 8'd211;  #10 
a = 8'd165; b = 8'd212;  #10 
a = 8'd165; b = 8'd213;  #10 
a = 8'd165; b = 8'd214;  #10 
a = 8'd165; b = 8'd215;  #10 
a = 8'd165; b = 8'd216;  #10 
a = 8'd165; b = 8'd217;  #10 
a = 8'd165; b = 8'd218;  #10 
a = 8'd165; b = 8'd219;  #10 
a = 8'd165; b = 8'd220;  #10 
a = 8'd165; b = 8'd221;  #10 
a = 8'd165; b = 8'd222;  #10 
a = 8'd165; b = 8'd223;  #10 
a = 8'd165; b = 8'd224;  #10 
a = 8'd165; b = 8'd225;  #10 
a = 8'd165; b = 8'd226;  #10 
a = 8'd165; b = 8'd227;  #10 
a = 8'd165; b = 8'd228;  #10 
a = 8'd165; b = 8'd229;  #10 
a = 8'd165; b = 8'd230;  #10 
a = 8'd165; b = 8'd231;  #10 
a = 8'd165; b = 8'd232;  #10 
a = 8'd165; b = 8'd233;  #10 
a = 8'd165; b = 8'd234;  #10 
a = 8'd165; b = 8'd235;  #10 
a = 8'd165; b = 8'd236;  #10 
a = 8'd165; b = 8'd237;  #10 
a = 8'd165; b = 8'd238;  #10 
a = 8'd165; b = 8'd239;  #10 
a = 8'd165; b = 8'd240;  #10 
a = 8'd165; b = 8'd241;  #10 
a = 8'd165; b = 8'd242;  #10 
a = 8'd165; b = 8'd243;  #10 
a = 8'd165; b = 8'd244;  #10 
a = 8'd165; b = 8'd245;  #10 
a = 8'd165; b = 8'd246;  #10 
a = 8'd165; b = 8'd247;  #10 
a = 8'd165; b = 8'd248;  #10 
a = 8'd165; b = 8'd249;  #10 
a = 8'd165; b = 8'd250;  #10 
a = 8'd165; b = 8'd251;  #10 
a = 8'd165; b = 8'd252;  #10 
a = 8'd165; b = 8'd253;  #10 
a = 8'd165; b = 8'd254;  #10 
a = 8'd165; b = 8'd255;  #10 
a = 8'd166; b = 8'd0;  #10 
a = 8'd166; b = 8'd1;  #10 
a = 8'd166; b = 8'd2;  #10 
a = 8'd166; b = 8'd3;  #10 
a = 8'd166; b = 8'd4;  #10 
a = 8'd166; b = 8'd5;  #10 
a = 8'd166; b = 8'd6;  #10 
a = 8'd166; b = 8'd7;  #10 
a = 8'd166; b = 8'd8;  #10 
a = 8'd166; b = 8'd9;  #10 
a = 8'd166; b = 8'd10;  #10 
a = 8'd166; b = 8'd11;  #10 
a = 8'd166; b = 8'd12;  #10 
a = 8'd166; b = 8'd13;  #10 
a = 8'd166; b = 8'd14;  #10 
a = 8'd166; b = 8'd15;  #10 
a = 8'd166; b = 8'd16;  #10 
a = 8'd166; b = 8'd17;  #10 
a = 8'd166; b = 8'd18;  #10 
a = 8'd166; b = 8'd19;  #10 
a = 8'd166; b = 8'd20;  #10 
a = 8'd166; b = 8'd21;  #10 
a = 8'd166; b = 8'd22;  #10 
a = 8'd166; b = 8'd23;  #10 
a = 8'd166; b = 8'd24;  #10 
a = 8'd166; b = 8'd25;  #10 
a = 8'd166; b = 8'd26;  #10 
a = 8'd166; b = 8'd27;  #10 
a = 8'd166; b = 8'd28;  #10 
a = 8'd166; b = 8'd29;  #10 
a = 8'd166; b = 8'd30;  #10 
a = 8'd166; b = 8'd31;  #10 
a = 8'd166; b = 8'd32;  #10 
a = 8'd166; b = 8'd33;  #10 
a = 8'd166; b = 8'd34;  #10 
a = 8'd166; b = 8'd35;  #10 
a = 8'd166; b = 8'd36;  #10 
a = 8'd166; b = 8'd37;  #10 
a = 8'd166; b = 8'd38;  #10 
a = 8'd166; b = 8'd39;  #10 
a = 8'd166; b = 8'd40;  #10 
a = 8'd166; b = 8'd41;  #10 
a = 8'd166; b = 8'd42;  #10 
a = 8'd166; b = 8'd43;  #10 
a = 8'd166; b = 8'd44;  #10 
a = 8'd166; b = 8'd45;  #10 
a = 8'd166; b = 8'd46;  #10 
a = 8'd166; b = 8'd47;  #10 
a = 8'd166; b = 8'd48;  #10 
a = 8'd166; b = 8'd49;  #10 
a = 8'd166; b = 8'd50;  #10 
a = 8'd166; b = 8'd51;  #10 
a = 8'd166; b = 8'd52;  #10 
a = 8'd166; b = 8'd53;  #10 
a = 8'd166; b = 8'd54;  #10 
a = 8'd166; b = 8'd55;  #10 
a = 8'd166; b = 8'd56;  #10 
a = 8'd166; b = 8'd57;  #10 
a = 8'd166; b = 8'd58;  #10 
a = 8'd166; b = 8'd59;  #10 
a = 8'd166; b = 8'd60;  #10 
a = 8'd166; b = 8'd61;  #10 
a = 8'd166; b = 8'd62;  #10 
a = 8'd166; b = 8'd63;  #10 
a = 8'd166; b = 8'd64;  #10 
a = 8'd166; b = 8'd65;  #10 
a = 8'd166; b = 8'd66;  #10 
a = 8'd166; b = 8'd67;  #10 
a = 8'd166; b = 8'd68;  #10 
a = 8'd166; b = 8'd69;  #10 
a = 8'd166; b = 8'd70;  #10 
a = 8'd166; b = 8'd71;  #10 
a = 8'd166; b = 8'd72;  #10 
a = 8'd166; b = 8'd73;  #10 
a = 8'd166; b = 8'd74;  #10 
a = 8'd166; b = 8'd75;  #10 
a = 8'd166; b = 8'd76;  #10 
a = 8'd166; b = 8'd77;  #10 
a = 8'd166; b = 8'd78;  #10 
a = 8'd166; b = 8'd79;  #10 
a = 8'd166; b = 8'd80;  #10 
a = 8'd166; b = 8'd81;  #10 
a = 8'd166; b = 8'd82;  #10 
a = 8'd166; b = 8'd83;  #10 
a = 8'd166; b = 8'd84;  #10 
a = 8'd166; b = 8'd85;  #10 
a = 8'd166; b = 8'd86;  #10 
a = 8'd166; b = 8'd87;  #10 
a = 8'd166; b = 8'd88;  #10 
a = 8'd166; b = 8'd89;  #10 
a = 8'd166; b = 8'd90;  #10 
a = 8'd166; b = 8'd91;  #10 
a = 8'd166; b = 8'd92;  #10 
a = 8'd166; b = 8'd93;  #10 
a = 8'd166; b = 8'd94;  #10 
a = 8'd166; b = 8'd95;  #10 
a = 8'd166; b = 8'd96;  #10 
a = 8'd166; b = 8'd97;  #10 
a = 8'd166; b = 8'd98;  #10 
a = 8'd166; b = 8'd99;  #10 
a = 8'd166; b = 8'd100;  #10 
a = 8'd166; b = 8'd101;  #10 
a = 8'd166; b = 8'd102;  #10 
a = 8'd166; b = 8'd103;  #10 
a = 8'd166; b = 8'd104;  #10 
a = 8'd166; b = 8'd105;  #10 
a = 8'd166; b = 8'd106;  #10 
a = 8'd166; b = 8'd107;  #10 
a = 8'd166; b = 8'd108;  #10 
a = 8'd166; b = 8'd109;  #10 
a = 8'd166; b = 8'd110;  #10 
a = 8'd166; b = 8'd111;  #10 
a = 8'd166; b = 8'd112;  #10 
a = 8'd166; b = 8'd113;  #10 
a = 8'd166; b = 8'd114;  #10 
a = 8'd166; b = 8'd115;  #10 
a = 8'd166; b = 8'd116;  #10 
a = 8'd166; b = 8'd117;  #10 
a = 8'd166; b = 8'd118;  #10 
a = 8'd166; b = 8'd119;  #10 
a = 8'd166; b = 8'd120;  #10 
a = 8'd166; b = 8'd121;  #10 
a = 8'd166; b = 8'd122;  #10 
a = 8'd166; b = 8'd123;  #10 
a = 8'd166; b = 8'd124;  #10 
a = 8'd166; b = 8'd125;  #10 
a = 8'd166; b = 8'd126;  #10 
a = 8'd166; b = 8'd127;  #10 
a = 8'd166; b = 8'd128;  #10 
a = 8'd166; b = 8'd129;  #10 
a = 8'd166; b = 8'd130;  #10 
a = 8'd166; b = 8'd131;  #10 
a = 8'd166; b = 8'd132;  #10 
a = 8'd166; b = 8'd133;  #10 
a = 8'd166; b = 8'd134;  #10 
a = 8'd166; b = 8'd135;  #10 
a = 8'd166; b = 8'd136;  #10 
a = 8'd166; b = 8'd137;  #10 
a = 8'd166; b = 8'd138;  #10 
a = 8'd166; b = 8'd139;  #10 
a = 8'd166; b = 8'd140;  #10 
a = 8'd166; b = 8'd141;  #10 
a = 8'd166; b = 8'd142;  #10 
a = 8'd166; b = 8'd143;  #10 
a = 8'd166; b = 8'd144;  #10 
a = 8'd166; b = 8'd145;  #10 
a = 8'd166; b = 8'd146;  #10 
a = 8'd166; b = 8'd147;  #10 
a = 8'd166; b = 8'd148;  #10 
a = 8'd166; b = 8'd149;  #10 
a = 8'd166; b = 8'd150;  #10 
a = 8'd166; b = 8'd151;  #10 
a = 8'd166; b = 8'd152;  #10 
a = 8'd166; b = 8'd153;  #10 
a = 8'd166; b = 8'd154;  #10 
a = 8'd166; b = 8'd155;  #10 
a = 8'd166; b = 8'd156;  #10 
a = 8'd166; b = 8'd157;  #10 
a = 8'd166; b = 8'd158;  #10 
a = 8'd166; b = 8'd159;  #10 
a = 8'd166; b = 8'd160;  #10 
a = 8'd166; b = 8'd161;  #10 
a = 8'd166; b = 8'd162;  #10 
a = 8'd166; b = 8'd163;  #10 
a = 8'd166; b = 8'd164;  #10 
a = 8'd166; b = 8'd165;  #10 
a = 8'd166; b = 8'd166;  #10 
a = 8'd166; b = 8'd167;  #10 
a = 8'd166; b = 8'd168;  #10 
a = 8'd166; b = 8'd169;  #10 
a = 8'd166; b = 8'd170;  #10 
a = 8'd166; b = 8'd171;  #10 
a = 8'd166; b = 8'd172;  #10 
a = 8'd166; b = 8'd173;  #10 
a = 8'd166; b = 8'd174;  #10 
a = 8'd166; b = 8'd175;  #10 
a = 8'd166; b = 8'd176;  #10 
a = 8'd166; b = 8'd177;  #10 
a = 8'd166; b = 8'd178;  #10 
a = 8'd166; b = 8'd179;  #10 
a = 8'd166; b = 8'd180;  #10 
a = 8'd166; b = 8'd181;  #10 
a = 8'd166; b = 8'd182;  #10 
a = 8'd166; b = 8'd183;  #10 
a = 8'd166; b = 8'd184;  #10 
a = 8'd166; b = 8'd185;  #10 
a = 8'd166; b = 8'd186;  #10 
a = 8'd166; b = 8'd187;  #10 
a = 8'd166; b = 8'd188;  #10 
a = 8'd166; b = 8'd189;  #10 
a = 8'd166; b = 8'd190;  #10 
a = 8'd166; b = 8'd191;  #10 
a = 8'd166; b = 8'd192;  #10 
a = 8'd166; b = 8'd193;  #10 
a = 8'd166; b = 8'd194;  #10 
a = 8'd166; b = 8'd195;  #10 
a = 8'd166; b = 8'd196;  #10 
a = 8'd166; b = 8'd197;  #10 
a = 8'd166; b = 8'd198;  #10 
a = 8'd166; b = 8'd199;  #10 
a = 8'd166; b = 8'd200;  #10 
a = 8'd166; b = 8'd201;  #10 
a = 8'd166; b = 8'd202;  #10 
a = 8'd166; b = 8'd203;  #10 
a = 8'd166; b = 8'd204;  #10 
a = 8'd166; b = 8'd205;  #10 
a = 8'd166; b = 8'd206;  #10 
a = 8'd166; b = 8'd207;  #10 
a = 8'd166; b = 8'd208;  #10 
a = 8'd166; b = 8'd209;  #10 
a = 8'd166; b = 8'd210;  #10 
a = 8'd166; b = 8'd211;  #10 
a = 8'd166; b = 8'd212;  #10 
a = 8'd166; b = 8'd213;  #10 
a = 8'd166; b = 8'd214;  #10 
a = 8'd166; b = 8'd215;  #10 
a = 8'd166; b = 8'd216;  #10 
a = 8'd166; b = 8'd217;  #10 
a = 8'd166; b = 8'd218;  #10 
a = 8'd166; b = 8'd219;  #10 
a = 8'd166; b = 8'd220;  #10 
a = 8'd166; b = 8'd221;  #10 
a = 8'd166; b = 8'd222;  #10 
a = 8'd166; b = 8'd223;  #10 
a = 8'd166; b = 8'd224;  #10 
a = 8'd166; b = 8'd225;  #10 
a = 8'd166; b = 8'd226;  #10 
a = 8'd166; b = 8'd227;  #10 
a = 8'd166; b = 8'd228;  #10 
a = 8'd166; b = 8'd229;  #10 
a = 8'd166; b = 8'd230;  #10 
a = 8'd166; b = 8'd231;  #10 
a = 8'd166; b = 8'd232;  #10 
a = 8'd166; b = 8'd233;  #10 
a = 8'd166; b = 8'd234;  #10 
a = 8'd166; b = 8'd235;  #10 
a = 8'd166; b = 8'd236;  #10 
a = 8'd166; b = 8'd237;  #10 
a = 8'd166; b = 8'd238;  #10 
a = 8'd166; b = 8'd239;  #10 
a = 8'd166; b = 8'd240;  #10 
a = 8'd166; b = 8'd241;  #10 
a = 8'd166; b = 8'd242;  #10 
a = 8'd166; b = 8'd243;  #10 
a = 8'd166; b = 8'd244;  #10 
a = 8'd166; b = 8'd245;  #10 
a = 8'd166; b = 8'd246;  #10 
a = 8'd166; b = 8'd247;  #10 
a = 8'd166; b = 8'd248;  #10 
a = 8'd166; b = 8'd249;  #10 
a = 8'd166; b = 8'd250;  #10 
a = 8'd166; b = 8'd251;  #10 
a = 8'd166; b = 8'd252;  #10 
a = 8'd166; b = 8'd253;  #10 
a = 8'd166; b = 8'd254;  #10 
a = 8'd166; b = 8'd255;  #10 
a = 8'd167; b = 8'd0;  #10 
a = 8'd167; b = 8'd1;  #10 
a = 8'd167; b = 8'd2;  #10 
a = 8'd167; b = 8'd3;  #10 
a = 8'd167; b = 8'd4;  #10 
a = 8'd167; b = 8'd5;  #10 
a = 8'd167; b = 8'd6;  #10 
a = 8'd167; b = 8'd7;  #10 
a = 8'd167; b = 8'd8;  #10 
a = 8'd167; b = 8'd9;  #10 
a = 8'd167; b = 8'd10;  #10 
a = 8'd167; b = 8'd11;  #10 
a = 8'd167; b = 8'd12;  #10 
a = 8'd167; b = 8'd13;  #10 
a = 8'd167; b = 8'd14;  #10 
a = 8'd167; b = 8'd15;  #10 
a = 8'd167; b = 8'd16;  #10 
a = 8'd167; b = 8'd17;  #10 
a = 8'd167; b = 8'd18;  #10 
a = 8'd167; b = 8'd19;  #10 
a = 8'd167; b = 8'd20;  #10 
a = 8'd167; b = 8'd21;  #10 
a = 8'd167; b = 8'd22;  #10 
a = 8'd167; b = 8'd23;  #10 
a = 8'd167; b = 8'd24;  #10 
a = 8'd167; b = 8'd25;  #10 
a = 8'd167; b = 8'd26;  #10 
a = 8'd167; b = 8'd27;  #10 
a = 8'd167; b = 8'd28;  #10 
a = 8'd167; b = 8'd29;  #10 
a = 8'd167; b = 8'd30;  #10 
a = 8'd167; b = 8'd31;  #10 
a = 8'd167; b = 8'd32;  #10 
a = 8'd167; b = 8'd33;  #10 
a = 8'd167; b = 8'd34;  #10 
a = 8'd167; b = 8'd35;  #10 
a = 8'd167; b = 8'd36;  #10 
a = 8'd167; b = 8'd37;  #10 
a = 8'd167; b = 8'd38;  #10 
a = 8'd167; b = 8'd39;  #10 
a = 8'd167; b = 8'd40;  #10 
a = 8'd167; b = 8'd41;  #10 
a = 8'd167; b = 8'd42;  #10 
a = 8'd167; b = 8'd43;  #10 
a = 8'd167; b = 8'd44;  #10 
a = 8'd167; b = 8'd45;  #10 
a = 8'd167; b = 8'd46;  #10 
a = 8'd167; b = 8'd47;  #10 
a = 8'd167; b = 8'd48;  #10 
a = 8'd167; b = 8'd49;  #10 
a = 8'd167; b = 8'd50;  #10 
a = 8'd167; b = 8'd51;  #10 
a = 8'd167; b = 8'd52;  #10 
a = 8'd167; b = 8'd53;  #10 
a = 8'd167; b = 8'd54;  #10 
a = 8'd167; b = 8'd55;  #10 
a = 8'd167; b = 8'd56;  #10 
a = 8'd167; b = 8'd57;  #10 
a = 8'd167; b = 8'd58;  #10 
a = 8'd167; b = 8'd59;  #10 
a = 8'd167; b = 8'd60;  #10 
a = 8'd167; b = 8'd61;  #10 
a = 8'd167; b = 8'd62;  #10 
a = 8'd167; b = 8'd63;  #10 
a = 8'd167; b = 8'd64;  #10 
a = 8'd167; b = 8'd65;  #10 
a = 8'd167; b = 8'd66;  #10 
a = 8'd167; b = 8'd67;  #10 
a = 8'd167; b = 8'd68;  #10 
a = 8'd167; b = 8'd69;  #10 
a = 8'd167; b = 8'd70;  #10 
a = 8'd167; b = 8'd71;  #10 
a = 8'd167; b = 8'd72;  #10 
a = 8'd167; b = 8'd73;  #10 
a = 8'd167; b = 8'd74;  #10 
a = 8'd167; b = 8'd75;  #10 
a = 8'd167; b = 8'd76;  #10 
a = 8'd167; b = 8'd77;  #10 
a = 8'd167; b = 8'd78;  #10 
a = 8'd167; b = 8'd79;  #10 
a = 8'd167; b = 8'd80;  #10 
a = 8'd167; b = 8'd81;  #10 
a = 8'd167; b = 8'd82;  #10 
a = 8'd167; b = 8'd83;  #10 
a = 8'd167; b = 8'd84;  #10 
a = 8'd167; b = 8'd85;  #10 
a = 8'd167; b = 8'd86;  #10 
a = 8'd167; b = 8'd87;  #10 
a = 8'd167; b = 8'd88;  #10 
a = 8'd167; b = 8'd89;  #10 
a = 8'd167; b = 8'd90;  #10 
a = 8'd167; b = 8'd91;  #10 
a = 8'd167; b = 8'd92;  #10 
a = 8'd167; b = 8'd93;  #10 
a = 8'd167; b = 8'd94;  #10 
a = 8'd167; b = 8'd95;  #10 
a = 8'd167; b = 8'd96;  #10 
a = 8'd167; b = 8'd97;  #10 
a = 8'd167; b = 8'd98;  #10 
a = 8'd167; b = 8'd99;  #10 
a = 8'd167; b = 8'd100;  #10 
a = 8'd167; b = 8'd101;  #10 
a = 8'd167; b = 8'd102;  #10 
a = 8'd167; b = 8'd103;  #10 
a = 8'd167; b = 8'd104;  #10 
a = 8'd167; b = 8'd105;  #10 
a = 8'd167; b = 8'd106;  #10 
a = 8'd167; b = 8'd107;  #10 
a = 8'd167; b = 8'd108;  #10 
a = 8'd167; b = 8'd109;  #10 
a = 8'd167; b = 8'd110;  #10 
a = 8'd167; b = 8'd111;  #10 
a = 8'd167; b = 8'd112;  #10 
a = 8'd167; b = 8'd113;  #10 
a = 8'd167; b = 8'd114;  #10 
a = 8'd167; b = 8'd115;  #10 
a = 8'd167; b = 8'd116;  #10 
a = 8'd167; b = 8'd117;  #10 
a = 8'd167; b = 8'd118;  #10 
a = 8'd167; b = 8'd119;  #10 
a = 8'd167; b = 8'd120;  #10 
a = 8'd167; b = 8'd121;  #10 
a = 8'd167; b = 8'd122;  #10 
a = 8'd167; b = 8'd123;  #10 
a = 8'd167; b = 8'd124;  #10 
a = 8'd167; b = 8'd125;  #10 
a = 8'd167; b = 8'd126;  #10 
a = 8'd167; b = 8'd127;  #10 
a = 8'd167; b = 8'd128;  #10 
a = 8'd167; b = 8'd129;  #10 
a = 8'd167; b = 8'd130;  #10 
a = 8'd167; b = 8'd131;  #10 
a = 8'd167; b = 8'd132;  #10 
a = 8'd167; b = 8'd133;  #10 
a = 8'd167; b = 8'd134;  #10 
a = 8'd167; b = 8'd135;  #10 
a = 8'd167; b = 8'd136;  #10 
a = 8'd167; b = 8'd137;  #10 
a = 8'd167; b = 8'd138;  #10 
a = 8'd167; b = 8'd139;  #10 
a = 8'd167; b = 8'd140;  #10 
a = 8'd167; b = 8'd141;  #10 
a = 8'd167; b = 8'd142;  #10 
a = 8'd167; b = 8'd143;  #10 
a = 8'd167; b = 8'd144;  #10 
a = 8'd167; b = 8'd145;  #10 
a = 8'd167; b = 8'd146;  #10 
a = 8'd167; b = 8'd147;  #10 
a = 8'd167; b = 8'd148;  #10 
a = 8'd167; b = 8'd149;  #10 
a = 8'd167; b = 8'd150;  #10 
a = 8'd167; b = 8'd151;  #10 
a = 8'd167; b = 8'd152;  #10 
a = 8'd167; b = 8'd153;  #10 
a = 8'd167; b = 8'd154;  #10 
a = 8'd167; b = 8'd155;  #10 
a = 8'd167; b = 8'd156;  #10 
a = 8'd167; b = 8'd157;  #10 
a = 8'd167; b = 8'd158;  #10 
a = 8'd167; b = 8'd159;  #10 
a = 8'd167; b = 8'd160;  #10 
a = 8'd167; b = 8'd161;  #10 
a = 8'd167; b = 8'd162;  #10 
a = 8'd167; b = 8'd163;  #10 
a = 8'd167; b = 8'd164;  #10 
a = 8'd167; b = 8'd165;  #10 
a = 8'd167; b = 8'd166;  #10 
a = 8'd167; b = 8'd167;  #10 
a = 8'd167; b = 8'd168;  #10 
a = 8'd167; b = 8'd169;  #10 
a = 8'd167; b = 8'd170;  #10 
a = 8'd167; b = 8'd171;  #10 
a = 8'd167; b = 8'd172;  #10 
a = 8'd167; b = 8'd173;  #10 
a = 8'd167; b = 8'd174;  #10 
a = 8'd167; b = 8'd175;  #10 
a = 8'd167; b = 8'd176;  #10 
a = 8'd167; b = 8'd177;  #10 
a = 8'd167; b = 8'd178;  #10 
a = 8'd167; b = 8'd179;  #10 
a = 8'd167; b = 8'd180;  #10 
a = 8'd167; b = 8'd181;  #10 
a = 8'd167; b = 8'd182;  #10 
a = 8'd167; b = 8'd183;  #10 
a = 8'd167; b = 8'd184;  #10 
a = 8'd167; b = 8'd185;  #10 
a = 8'd167; b = 8'd186;  #10 
a = 8'd167; b = 8'd187;  #10 
a = 8'd167; b = 8'd188;  #10 
a = 8'd167; b = 8'd189;  #10 
a = 8'd167; b = 8'd190;  #10 
a = 8'd167; b = 8'd191;  #10 
a = 8'd167; b = 8'd192;  #10 
a = 8'd167; b = 8'd193;  #10 
a = 8'd167; b = 8'd194;  #10 
a = 8'd167; b = 8'd195;  #10 
a = 8'd167; b = 8'd196;  #10 
a = 8'd167; b = 8'd197;  #10 
a = 8'd167; b = 8'd198;  #10 
a = 8'd167; b = 8'd199;  #10 
a = 8'd167; b = 8'd200;  #10 
a = 8'd167; b = 8'd201;  #10 
a = 8'd167; b = 8'd202;  #10 
a = 8'd167; b = 8'd203;  #10 
a = 8'd167; b = 8'd204;  #10 
a = 8'd167; b = 8'd205;  #10 
a = 8'd167; b = 8'd206;  #10 
a = 8'd167; b = 8'd207;  #10 
a = 8'd167; b = 8'd208;  #10 
a = 8'd167; b = 8'd209;  #10 
a = 8'd167; b = 8'd210;  #10 
a = 8'd167; b = 8'd211;  #10 
a = 8'd167; b = 8'd212;  #10 
a = 8'd167; b = 8'd213;  #10 
a = 8'd167; b = 8'd214;  #10 
a = 8'd167; b = 8'd215;  #10 
a = 8'd167; b = 8'd216;  #10 
a = 8'd167; b = 8'd217;  #10 
a = 8'd167; b = 8'd218;  #10 
a = 8'd167; b = 8'd219;  #10 
a = 8'd167; b = 8'd220;  #10 
a = 8'd167; b = 8'd221;  #10 
a = 8'd167; b = 8'd222;  #10 
a = 8'd167; b = 8'd223;  #10 
a = 8'd167; b = 8'd224;  #10 
a = 8'd167; b = 8'd225;  #10 
a = 8'd167; b = 8'd226;  #10 
a = 8'd167; b = 8'd227;  #10 
a = 8'd167; b = 8'd228;  #10 
a = 8'd167; b = 8'd229;  #10 
a = 8'd167; b = 8'd230;  #10 
a = 8'd167; b = 8'd231;  #10 
a = 8'd167; b = 8'd232;  #10 
a = 8'd167; b = 8'd233;  #10 
a = 8'd167; b = 8'd234;  #10 
a = 8'd167; b = 8'd235;  #10 
a = 8'd167; b = 8'd236;  #10 
a = 8'd167; b = 8'd237;  #10 
a = 8'd167; b = 8'd238;  #10 
a = 8'd167; b = 8'd239;  #10 
a = 8'd167; b = 8'd240;  #10 
a = 8'd167; b = 8'd241;  #10 
a = 8'd167; b = 8'd242;  #10 
a = 8'd167; b = 8'd243;  #10 
a = 8'd167; b = 8'd244;  #10 
a = 8'd167; b = 8'd245;  #10 
a = 8'd167; b = 8'd246;  #10 
a = 8'd167; b = 8'd247;  #10 
a = 8'd167; b = 8'd248;  #10 
a = 8'd167; b = 8'd249;  #10 
a = 8'd167; b = 8'd250;  #10 
a = 8'd167; b = 8'd251;  #10 
a = 8'd167; b = 8'd252;  #10 
a = 8'd167; b = 8'd253;  #10 
a = 8'd167; b = 8'd254;  #10 
a = 8'd167; b = 8'd255;  #10 
a = 8'd168; b = 8'd0;  #10 
a = 8'd168; b = 8'd1;  #10 
a = 8'd168; b = 8'd2;  #10 
a = 8'd168; b = 8'd3;  #10 
a = 8'd168; b = 8'd4;  #10 
a = 8'd168; b = 8'd5;  #10 
a = 8'd168; b = 8'd6;  #10 
a = 8'd168; b = 8'd7;  #10 
a = 8'd168; b = 8'd8;  #10 
a = 8'd168; b = 8'd9;  #10 
a = 8'd168; b = 8'd10;  #10 
a = 8'd168; b = 8'd11;  #10 
a = 8'd168; b = 8'd12;  #10 
a = 8'd168; b = 8'd13;  #10 
a = 8'd168; b = 8'd14;  #10 
a = 8'd168; b = 8'd15;  #10 
a = 8'd168; b = 8'd16;  #10 
a = 8'd168; b = 8'd17;  #10 
a = 8'd168; b = 8'd18;  #10 
a = 8'd168; b = 8'd19;  #10 
a = 8'd168; b = 8'd20;  #10 
a = 8'd168; b = 8'd21;  #10 
a = 8'd168; b = 8'd22;  #10 
a = 8'd168; b = 8'd23;  #10 
a = 8'd168; b = 8'd24;  #10 
a = 8'd168; b = 8'd25;  #10 
a = 8'd168; b = 8'd26;  #10 
a = 8'd168; b = 8'd27;  #10 
a = 8'd168; b = 8'd28;  #10 
a = 8'd168; b = 8'd29;  #10 
a = 8'd168; b = 8'd30;  #10 
a = 8'd168; b = 8'd31;  #10 
a = 8'd168; b = 8'd32;  #10 
a = 8'd168; b = 8'd33;  #10 
a = 8'd168; b = 8'd34;  #10 
a = 8'd168; b = 8'd35;  #10 
a = 8'd168; b = 8'd36;  #10 
a = 8'd168; b = 8'd37;  #10 
a = 8'd168; b = 8'd38;  #10 
a = 8'd168; b = 8'd39;  #10 
a = 8'd168; b = 8'd40;  #10 
a = 8'd168; b = 8'd41;  #10 
a = 8'd168; b = 8'd42;  #10 
a = 8'd168; b = 8'd43;  #10 
a = 8'd168; b = 8'd44;  #10 
a = 8'd168; b = 8'd45;  #10 
a = 8'd168; b = 8'd46;  #10 
a = 8'd168; b = 8'd47;  #10 
a = 8'd168; b = 8'd48;  #10 
a = 8'd168; b = 8'd49;  #10 
a = 8'd168; b = 8'd50;  #10 
a = 8'd168; b = 8'd51;  #10 
a = 8'd168; b = 8'd52;  #10 
a = 8'd168; b = 8'd53;  #10 
a = 8'd168; b = 8'd54;  #10 
a = 8'd168; b = 8'd55;  #10 
a = 8'd168; b = 8'd56;  #10 
a = 8'd168; b = 8'd57;  #10 
a = 8'd168; b = 8'd58;  #10 
a = 8'd168; b = 8'd59;  #10 
a = 8'd168; b = 8'd60;  #10 
a = 8'd168; b = 8'd61;  #10 
a = 8'd168; b = 8'd62;  #10 
a = 8'd168; b = 8'd63;  #10 
a = 8'd168; b = 8'd64;  #10 
a = 8'd168; b = 8'd65;  #10 
a = 8'd168; b = 8'd66;  #10 
a = 8'd168; b = 8'd67;  #10 
a = 8'd168; b = 8'd68;  #10 
a = 8'd168; b = 8'd69;  #10 
a = 8'd168; b = 8'd70;  #10 
a = 8'd168; b = 8'd71;  #10 
a = 8'd168; b = 8'd72;  #10 
a = 8'd168; b = 8'd73;  #10 
a = 8'd168; b = 8'd74;  #10 
a = 8'd168; b = 8'd75;  #10 
a = 8'd168; b = 8'd76;  #10 
a = 8'd168; b = 8'd77;  #10 
a = 8'd168; b = 8'd78;  #10 
a = 8'd168; b = 8'd79;  #10 
a = 8'd168; b = 8'd80;  #10 
a = 8'd168; b = 8'd81;  #10 
a = 8'd168; b = 8'd82;  #10 
a = 8'd168; b = 8'd83;  #10 
a = 8'd168; b = 8'd84;  #10 
a = 8'd168; b = 8'd85;  #10 
a = 8'd168; b = 8'd86;  #10 
a = 8'd168; b = 8'd87;  #10 
a = 8'd168; b = 8'd88;  #10 
a = 8'd168; b = 8'd89;  #10 
a = 8'd168; b = 8'd90;  #10 
a = 8'd168; b = 8'd91;  #10 
a = 8'd168; b = 8'd92;  #10 
a = 8'd168; b = 8'd93;  #10 
a = 8'd168; b = 8'd94;  #10 
a = 8'd168; b = 8'd95;  #10 
a = 8'd168; b = 8'd96;  #10 
a = 8'd168; b = 8'd97;  #10 
a = 8'd168; b = 8'd98;  #10 
a = 8'd168; b = 8'd99;  #10 
a = 8'd168; b = 8'd100;  #10 
a = 8'd168; b = 8'd101;  #10 
a = 8'd168; b = 8'd102;  #10 
a = 8'd168; b = 8'd103;  #10 
a = 8'd168; b = 8'd104;  #10 
a = 8'd168; b = 8'd105;  #10 
a = 8'd168; b = 8'd106;  #10 
a = 8'd168; b = 8'd107;  #10 
a = 8'd168; b = 8'd108;  #10 
a = 8'd168; b = 8'd109;  #10 
a = 8'd168; b = 8'd110;  #10 
a = 8'd168; b = 8'd111;  #10 
a = 8'd168; b = 8'd112;  #10 
a = 8'd168; b = 8'd113;  #10 
a = 8'd168; b = 8'd114;  #10 
a = 8'd168; b = 8'd115;  #10 
a = 8'd168; b = 8'd116;  #10 
a = 8'd168; b = 8'd117;  #10 
a = 8'd168; b = 8'd118;  #10 
a = 8'd168; b = 8'd119;  #10 
a = 8'd168; b = 8'd120;  #10 
a = 8'd168; b = 8'd121;  #10 
a = 8'd168; b = 8'd122;  #10 
a = 8'd168; b = 8'd123;  #10 
a = 8'd168; b = 8'd124;  #10 
a = 8'd168; b = 8'd125;  #10 
a = 8'd168; b = 8'd126;  #10 
a = 8'd168; b = 8'd127;  #10 
a = 8'd168; b = 8'd128;  #10 
a = 8'd168; b = 8'd129;  #10 
a = 8'd168; b = 8'd130;  #10 
a = 8'd168; b = 8'd131;  #10 
a = 8'd168; b = 8'd132;  #10 
a = 8'd168; b = 8'd133;  #10 
a = 8'd168; b = 8'd134;  #10 
a = 8'd168; b = 8'd135;  #10 
a = 8'd168; b = 8'd136;  #10 
a = 8'd168; b = 8'd137;  #10 
a = 8'd168; b = 8'd138;  #10 
a = 8'd168; b = 8'd139;  #10 
a = 8'd168; b = 8'd140;  #10 
a = 8'd168; b = 8'd141;  #10 
a = 8'd168; b = 8'd142;  #10 
a = 8'd168; b = 8'd143;  #10 
a = 8'd168; b = 8'd144;  #10 
a = 8'd168; b = 8'd145;  #10 
a = 8'd168; b = 8'd146;  #10 
a = 8'd168; b = 8'd147;  #10 
a = 8'd168; b = 8'd148;  #10 
a = 8'd168; b = 8'd149;  #10 
a = 8'd168; b = 8'd150;  #10 
a = 8'd168; b = 8'd151;  #10 
a = 8'd168; b = 8'd152;  #10 
a = 8'd168; b = 8'd153;  #10 
a = 8'd168; b = 8'd154;  #10 
a = 8'd168; b = 8'd155;  #10 
a = 8'd168; b = 8'd156;  #10 
a = 8'd168; b = 8'd157;  #10 
a = 8'd168; b = 8'd158;  #10 
a = 8'd168; b = 8'd159;  #10 
a = 8'd168; b = 8'd160;  #10 
a = 8'd168; b = 8'd161;  #10 
a = 8'd168; b = 8'd162;  #10 
a = 8'd168; b = 8'd163;  #10 
a = 8'd168; b = 8'd164;  #10 
a = 8'd168; b = 8'd165;  #10 
a = 8'd168; b = 8'd166;  #10 
a = 8'd168; b = 8'd167;  #10 
a = 8'd168; b = 8'd168;  #10 
a = 8'd168; b = 8'd169;  #10 
a = 8'd168; b = 8'd170;  #10 
a = 8'd168; b = 8'd171;  #10 
a = 8'd168; b = 8'd172;  #10 
a = 8'd168; b = 8'd173;  #10 
a = 8'd168; b = 8'd174;  #10 
a = 8'd168; b = 8'd175;  #10 
a = 8'd168; b = 8'd176;  #10 
a = 8'd168; b = 8'd177;  #10 
a = 8'd168; b = 8'd178;  #10 
a = 8'd168; b = 8'd179;  #10 
a = 8'd168; b = 8'd180;  #10 
a = 8'd168; b = 8'd181;  #10 
a = 8'd168; b = 8'd182;  #10 
a = 8'd168; b = 8'd183;  #10 
a = 8'd168; b = 8'd184;  #10 
a = 8'd168; b = 8'd185;  #10 
a = 8'd168; b = 8'd186;  #10 
a = 8'd168; b = 8'd187;  #10 
a = 8'd168; b = 8'd188;  #10 
a = 8'd168; b = 8'd189;  #10 
a = 8'd168; b = 8'd190;  #10 
a = 8'd168; b = 8'd191;  #10 
a = 8'd168; b = 8'd192;  #10 
a = 8'd168; b = 8'd193;  #10 
a = 8'd168; b = 8'd194;  #10 
a = 8'd168; b = 8'd195;  #10 
a = 8'd168; b = 8'd196;  #10 
a = 8'd168; b = 8'd197;  #10 
a = 8'd168; b = 8'd198;  #10 
a = 8'd168; b = 8'd199;  #10 
a = 8'd168; b = 8'd200;  #10 
a = 8'd168; b = 8'd201;  #10 
a = 8'd168; b = 8'd202;  #10 
a = 8'd168; b = 8'd203;  #10 
a = 8'd168; b = 8'd204;  #10 
a = 8'd168; b = 8'd205;  #10 
a = 8'd168; b = 8'd206;  #10 
a = 8'd168; b = 8'd207;  #10 
a = 8'd168; b = 8'd208;  #10 
a = 8'd168; b = 8'd209;  #10 
a = 8'd168; b = 8'd210;  #10 
a = 8'd168; b = 8'd211;  #10 
a = 8'd168; b = 8'd212;  #10 
a = 8'd168; b = 8'd213;  #10 
a = 8'd168; b = 8'd214;  #10 
a = 8'd168; b = 8'd215;  #10 
a = 8'd168; b = 8'd216;  #10 
a = 8'd168; b = 8'd217;  #10 
a = 8'd168; b = 8'd218;  #10 
a = 8'd168; b = 8'd219;  #10 
a = 8'd168; b = 8'd220;  #10 
a = 8'd168; b = 8'd221;  #10 
a = 8'd168; b = 8'd222;  #10 
a = 8'd168; b = 8'd223;  #10 
a = 8'd168; b = 8'd224;  #10 
a = 8'd168; b = 8'd225;  #10 
a = 8'd168; b = 8'd226;  #10 
a = 8'd168; b = 8'd227;  #10 
a = 8'd168; b = 8'd228;  #10 
a = 8'd168; b = 8'd229;  #10 
a = 8'd168; b = 8'd230;  #10 
a = 8'd168; b = 8'd231;  #10 
a = 8'd168; b = 8'd232;  #10 
a = 8'd168; b = 8'd233;  #10 
a = 8'd168; b = 8'd234;  #10 
a = 8'd168; b = 8'd235;  #10 
a = 8'd168; b = 8'd236;  #10 
a = 8'd168; b = 8'd237;  #10 
a = 8'd168; b = 8'd238;  #10 
a = 8'd168; b = 8'd239;  #10 
a = 8'd168; b = 8'd240;  #10 
a = 8'd168; b = 8'd241;  #10 
a = 8'd168; b = 8'd242;  #10 
a = 8'd168; b = 8'd243;  #10 
a = 8'd168; b = 8'd244;  #10 
a = 8'd168; b = 8'd245;  #10 
a = 8'd168; b = 8'd246;  #10 
a = 8'd168; b = 8'd247;  #10 
a = 8'd168; b = 8'd248;  #10 
a = 8'd168; b = 8'd249;  #10 
a = 8'd168; b = 8'd250;  #10 
a = 8'd168; b = 8'd251;  #10 
a = 8'd168; b = 8'd252;  #10 
a = 8'd168; b = 8'd253;  #10 
a = 8'd168; b = 8'd254;  #10 
a = 8'd168; b = 8'd255;  #10 
a = 8'd169; b = 8'd0;  #10 
a = 8'd169; b = 8'd1;  #10 
a = 8'd169; b = 8'd2;  #10 
a = 8'd169; b = 8'd3;  #10 
a = 8'd169; b = 8'd4;  #10 
a = 8'd169; b = 8'd5;  #10 
a = 8'd169; b = 8'd6;  #10 
a = 8'd169; b = 8'd7;  #10 
a = 8'd169; b = 8'd8;  #10 
a = 8'd169; b = 8'd9;  #10 
a = 8'd169; b = 8'd10;  #10 
a = 8'd169; b = 8'd11;  #10 
a = 8'd169; b = 8'd12;  #10 
a = 8'd169; b = 8'd13;  #10 
a = 8'd169; b = 8'd14;  #10 
a = 8'd169; b = 8'd15;  #10 
a = 8'd169; b = 8'd16;  #10 
a = 8'd169; b = 8'd17;  #10 
a = 8'd169; b = 8'd18;  #10 
a = 8'd169; b = 8'd19;  #10 
a = 8'd169; b = 8'd20;  #10 
a = 8'd169; b = 8'd21;  #10 
a = 8'd169; b = 8'd22;  #10 
a = 8'd169; b = 8'd23;  #10 
a = 8'd169; b = 8'd24;  #10 
a = 8'd169; b = 8'd25;  #10 
a = 8'd169; b = 8'd26;  #10 
a = 8'd169; b = 8'd27;  #10 
a = 8'd169; b = 8'd28;  #10 
a = 8'd169; b = 8'd29;  #10 
a = 8'd169; b = 8'd30;  #10 
a = 8'd169; b = 8'd31;  #10 
a = 8'd169; b = 8'd32;  #10 
a = 8'd169; b = 8'd33;  #10 
a = 8'd169; b = 8'd34;  #10 
a = 8'd169; b = 8'd35;  #10 
a = 8'd169; b = 8'd36;  #10 
a = 8'd169; b = 8'd37;  #10 
a = 8'd169; b = 8'd38;  #10 
a = 8'd169; b = 8'd39;  #10 
a = 8'd169; b = 8'd40;  #10 
a = 8'd169; b = 8'd41;  #10 
a = 8'd169; b = 8'd42;  #10 
a = 8'd169; b = 8'd43;  #10 
a = 8'd169; b = 8'd44;  #10 
a = 8'd169; b = 8'd45;  #10 
a = 8'd169; b = 8'd46;  #10 
a = 8'd169; b = 8'd47;  #10 
a = 8'd169; b = 8'd48;  #10 
a = 8'd169; b = 8'd49;  #10 
a = 8'd169; b = 8'd50;  #10 
a = 8'd169; b = 8'd51;  #10 
a = 8'd169; b = 8'd52;  #10 
a = 8'd169; b = 8'd53;  #10 
a = 8'd169; b = 8'd54;  #10 
a = 8'd169; b = 8'd55;  #10 
a = 8'd169; b = 8'd56;  #10 
a = 8'd169; b = 8'd57;  #10 
a = 8'd169; b = 8'd58;  #10 
a = 8'd169; b = 8'd59;  #10 
a = 8'd169; b = 8'd60;  #10 
a = 8'd169; b = 8'd61;  #10 
a = 8'd169; b = 8'd62;  #10 
a = 8'd169; b = 8'd63;  #10 
a = 8'd169; b = 8'd64;  #10 
a = 8'd169; b = 8'd65;  #10 
a = 8'd169; b = 8'd66;  #10 
a = 8'd169; b = 8'd67;  #10 
a = 8'd169; b = 8'd68;  #10 
a = 8'd169; b = 8'd69;  #10 
a = 8'd169; b = 8'd70;  #10 
a = 8'd169; b = 8'd71;  #10 
a = 8'd169; b = 8'd72;  #10 
a = 8'd169; b = 8'd73;  #10 
a = 8'd169; b = 8'd74;  #10 
a = 8'd169; b = 8'd75;  #10 
a = 8'd169; b = 8'd76;  #10 
a = 8'd169; b = 8'd77;  #10 
a = 8'd169; b = 8'd78;  #10 
a = 8'd169; b = 8'd79;  #10 
a = 8'd169; b = 8'd80;  #10 
a = 8'd169; b = 8'd81;  #10 
a = 8'd169; b = 8'd82;  #10 
a = 8'd169; b = 8'd83;  #10 
a = 8'd169; b = 8'd84;  #10 
a = 8'd169; b = 8'd85;  #10 
a = 8'd169; b = 8'd86;  #10 
a = 8'd169; b = 8'd87;  #10 
a = 8'd169; b = 8'd88;  #10 
a = 8'd169; b = 8'd89;  #10 
a = 8'd169; b = 8'd90;  #10 
a = 8'd169; b = 8'd91;  #10 
a = 8'd169; b = 8'd92;  #10 
a = 8'd169; b = 8'd93;  #10 
a = 8'd169; b = 8'd94;  #10 
a = 8'd169; b = 8'd95;  #10 
a = 8'd169; b = 8'd96;  #10 
a = 8'd169; b = 8'd97;  #10 
a = 8'd169; b = 8'd98;  #10 
a = 8'd169; b = 8'd99;  #10 
a = 8'd169; b = 8'd100;  #10 
a = 8'd169; b = 8'd101;  #10 
a = 8'd169; b = 8'd102;  #10 
a = 8'd169; b = 8'd103;  #10 
a = 8'd169; b = 8'd104;  #10 
a = 8'd169; b = 8'd105;  #10 
a = 8'd169; b = 8'd106;  #10 
a = 8'd169; b = 8'd107;  #10 
a = 8'd169; b = 8'd108;  #10 
a = 8'd169; b = 8'd109;  #10 
a = 8'd169; b = 8'd110;  #10 
a = 8'd169; b = 8'd111;  #10 
a = 8'd169; b = 8'd112;  #10 
a = 8'd169; b = 8'd113;  #10 
a = 8'd169; b = 8'd114;  #10 
a = 8'd169; b = 8'd115;  #10 
a = 8'd169; b = 8'd116;  #10 
a = 8'd169; b = 8'd117;  #10 
a = 8'd169; b = 8'd118;  #10 
a = 8'd169; b = 8'd119;  #10 
a = 8'd169; b = 8'd120;  #10 
a = 8'd169; b = 8'd121;  #10 
a = 8'd169; b = 8'd122;  #10 
a = 8'd169; b = 8'd123;  #10 
a = 8'd169; b = 8'd124;  #10 
a = 8'd169; b = 8'd125;  #10 
a = 8'd169; b = 8'd126;  #10 
a = 8'd169; b = 8'd127;  #10 
a = 8'd169; b = 8'd128;  #10 
a = 8'd169; b = 8'd129;  #10 
a = 8'd169; b = 8'd130;  #10 
a = 8'd169; b = 8'd131;  #10 
a = 8'd169; b = 8'd132;  #10 
a = 8'd169; b = 8'd133;  #10 
a = 8'd169; b = 8'd134;  #10 
a = 8'd169; b = 8'd135;  #10 
a = 8'd169; b = 8'd136;  #10 
a = 8'd169; b = 8'd137;  #10 
a = 8'd169; b = 8'd138;  #10 
a = 8'd169; b = 8'd139;  #10 
a = 8'd169; b = 8'd140;  #10 
a = 8'd169; b = 8'd141;  #10 
a = 8'd169; b = 8'd142;  #10 
a = 8'd169; b = 8'd143;  #10 
a = 8'd169; b = 8'd144;  #10 
a = 8'd169; b = 8'd145;  #10 
a = 8'd169; b = 8'd146;  #10 
a = 8'd169; b = 8'd147;  #10 
a = 8'd169; b = 8'd148;  #10 
a = 8'd169; b = 8'd149;  #10 
a = 8'd169; b = 8'd150;  #10 
a = 8'd169; b = 8'd151;  #10 
a = 8'd169; b = 8'd152;  #10 
a = 8'd169; b = 8'd153;  #10 
a = 8'd169; b = 8'd154;  #10 
a = 8'd169; b = 8'd155;  #10 
a = 8'd169; b = 8'd156;  #10 
a = 8'd169; b = 8'd157;  #10 
a = 8'd169; b = 8'd158;  #10 
a = 8'd169; b = 8'd159;  #10 
a = 8'd169; b = 8'd160;  #10 
a = 8'd169; b = 8'd161;  #10 
a = 8'd169; b = 8'd162;  #10 
a = 8'd169; b = 8'd163;  #10 
a = 8'd169; b = 8'd164;  #10 
a = 8'd169; b = 8'd165;  #10 
a = 8'd169; b = 8'd166;  #10 
a = 8'd169; b = 8'd167;  #10 
a = 8'd169; b = 8'd168;  #10 
a = 8'd169; b = 8'd169;  #10 
a = 8'd169; b = 8'd170;  #10 
a = 8'd169; b = 8'd171;  #10 
a = 8'd169; b = 8'd172;  #10 
a = 8'd169; b = 8'd173;  #10 
a = 8'd169; b = 8'd174;  #10 
a = 8'd169; b = 8'd175;  #10 
a = 8'd169; b = 8'd176;  #10 
a = 8'd169; b = 8'd177;  #10 
a = 8'd169; b = 8'd178;  #10 
a = 8'd169; b = 8'd179;  #10 
a = 8'd169; b = 8'd180;  #10 
a = 8'd169; b = 8'd181;  #10 
a = 8'd169; b = 8'd182;  #10 
a = 8'd169; b = 8'd183;  #10 
a = 8'd169; b = 8'd184;  #10 
a = 8'd169; b = 8'd185;  #10 
a = 8'd169; b = 8'd186;  #10 
a = 8'd169; b = 8'd187;  #10 
a = 8'd169; b = 8'd188;  #10 
a = 8'd169; b = 8'd189;  #10 
a = 8'd169; b = 8'd190;  #10 
a = 8'd169; b = 8'd191;  #10 
a = 8'd169; b = 8'd192;  #10 
a = 8'd169; b = 8'd193;  #10 
a = 8'd169; b = 8'd194;  #10 
a = 8'd169; b = 8'd195;  #10 
a = 8'd169; b = 8'd196;  #10 
a = 8'd169; b = 8'd197;  #10 
a = 8'd169; b = 8'd198;  #10 
a = 8'd169; b = 8'd199;  #10 
a = 8'd169; b = 8'd200;  #10 
a = 8'd169; b = 8'd201;  #10 
a = 8'd169; b = 8'd202;  #10 
a = 8'd169; b = 8'd203;  #10 
a = 8'd169; b = 8'd204;  #10 
a = 8'd169; b = 8'd205;  #10 
a = 8'd169; b = 8'd206;  #10 
a = 8'd169; b = 8'd207;  #10 
a = 8'd169; b = 8'd208;  #10 
a = 8'd169; b = 8'd209;  #10 
a = 8'd169; b = 8'd210;  #10 
a = 8'd169; b = 8'd211;  #10 
a = 8'd169; b = 8'd212;  #10 
a = 8'd169; b = 8'd213;  #10 
a = 8'd169; b = 8'd214;  #10 
a = 8'd169; b = 8'd215;  #10 
a = 8'd169; b = 8'd216;  #10 
a = 8'd169; b = 8'd217;  #10 
a = 8'd169; b = 8'd218;  #10 
a = 8'd169; b = 8'd219;  #10 
a = 8'd169; b = 8'd220;  #10 
a = 8'd169; b = 8'd221;  #10 
a = 8'd169; b = 8'd222;  #10 
a = 8'd169; b = 8'd223;  #10 
a = 8'd169; b = 8'd224;  #10 
a = 8'd169; b = 8'd225;  #10 
a = 8'd169; b = 8'd226;  #10 
a = 8'd169; b = 8'd227;  #10 
a = 8'd169; b = 8'd228;  #10 
a = 8'd169; b = 8'd229;  #10 
a = 8'd169; b = 8'd230;  #10 
a = 8'd169; b = 8'd231;  #10 
a = 8'd169; b = 8'd232;  #10 
a = 8'd169; b = 8'd233;  #10 
a = 8'd169; b = 8'd234;  #10 
a = 8'd169; b = 8'd235;  #10 
a = 8'd169; b = 8'd236;  #10 
a = 8'd169; b = 8'd237;  #10 
a = 8'd169; b = 8'd238;  #10 
a = 8'd169; b = 8'd239;  #10 
a = 8'd169; b = 8'd240;  #10 
a = 8'd169; b = 8'd241;  #10 
a = 8'd169; b = 8'd242;  #10 
a = 8'd169; b = 8'd243;  #10 
a = 8'd169; b = 8'd244;  #10 
a = 8'd169; b = 8'd245;  #10 
a = 8'd169; b = 8'd246;  #10 
a = 8'd169; b = 8'd247;  #10 
a = 8'd169; b = 8'd248;  #10 
a = 8'd169; b = 8'd249;  #10 
a = 8'd169; b = 8'd250;  #10 
a = 8'd169; b = 8'd251;  #10 
a = 8'd169; b = 8'd252;  #10 
a = 8'd169; b = 8'd253;  #10 
a = 8'd169; b = 8'd254;  #10 
a = 8'd169; b = 8'd255;  #10 
a = 8'd170; b = 8'd0;  #10 
a = 8'd170; b = 8'd1;  #10 
a = 8'd170; b = 8'd2;  #10 
a = 8'd170; b = 8'd3;  #10 
a = 8'd170; b = 8'd4;  #10 
a = 8'd170; b = 8'd5;  #10 
a = 8'd170; b = 8'd6;  #10 
a = 8'd170; b = 8'd7;  #10 
a = 8'd170; b = 8'd8;  #10 
a = 8'd170; b = 8'd9;  #10 
a = 8'd170; b = 8'd10;  #10 
a = 8'd170; b = 8'd11;  #10 
a = 8'd170; b = 8'd12;  #10 
a = 8'd170; b = 8'd13;  #10 
a = 8'd170; b = 8'd14;  #10 
a = 8'd170; b = 8'd15;  #10 
a = 8'd170; b = 8'd16;  #10 
a = 8'd170; b = 8'd17;  #10 
a = 8'd170; b = 8'd18;  #10 
a = 8'd170; b = 8'd19;  #10 
a = 8'd170; b = 8'd20;  #10 
a = 8'd170; b = 8'd21;  #10 
a = 8'd170; b = 8'd22;  #10 
a = 8'd170; b = 8'd23;  #10 
a = 8'd170; b = 8'd24;  #10 
a = 8'd170; b = 8'd25;  #10 
a = 8'd170; b = 8'd26;  #10 
a = 8'd170; b = 8'd27;  #10 
a = 8'd170; b = 8'd28;  #10 
a = 8'd170; b = 8'd29;  #10 
a = 8'd170; b = 8'd30;  #10 
a = 8'd170; b = 8'd31;  #10 
a = 8'd170; b = 8'd32;  #10 
a = 8'd170; b = 8'd33;  #10 
a = 8'd170; b = 8'd34;  #10 
a = 8'd170; b = 8'd35;  #10 
a = 8'd170; b = 8'd36;  #10 
a = 8'd170; b = 8'd37;  #10 
a = 8'd170; b = 8'd38;  #10 
a = 8'd170; b = 8'd39;  #10 
a = 8'd170; b = 8'd40;  #10 
a = 8'd170; b = 8'd41;  #10 
a = 8'd170; b = 8'd42;  #10 
a = 8'd170; b = 8'd43;  #10 
a = 8'd170; b = 8'd44;  #10 
a = 8'd170; b = 8'd45;  #10 
a = 8'd170; b = 8'd46;  #10 
a = 8'd170; b = 8'd47;  #10 
a = 8'd170; b = 8'd48;  #10 
a = 8'd170; b = 8'd49;  #10 
a = 8'd170; b = 8'd50;  #10 
a = 8'd170; b = 8'd51;  #10 
a = 8'd170; b = 8'd52;  #10 
a = 8'd170; b = 8'd53;  #10 
a = 8'd170; b = 8'd54;  #10 
a = 8'd170; b = 8'd55;  #10 
a = 8'd170; b = 8'd56;  #10 
a = 8'd170; b = 8'd57;  #10 
a = 8'd170; b = 8'd58;  #10 
a = 8'd170; b = 8'd59;  #10 
a = 8'd170; b = 8'd60;  #10 
a = 8'd170; b = 8'd61;  #10 
a = 8'd170; b = 8'd62;  #10 
a = 8'd170; b = 8'd63;  #10 
a = 8'd170; b = 8'd64;  #10 
a = 8'd170; b = 8'd65;  #10 
a = 8'd170; b = 8'd66;  #10 
a = 8'd170; b = 8'd67;  #10 
a = 8'd170; b = 8'd68;  #10 
a = 8'd170; b = 8'd69;  #10 
a = 8'd170; b = 8'd70;  #10 
a = 8'd170; b = 8'd71;  #10 
a = 8'd170; b = 8'd72;  #10 
a = 8'd170; b = 8'd73;  #10 
a = 8'd170; b = 8'd74;  #10 
a = 8'd170; b = 8'd75;  #10 
a = 8'd170; b = 8'd76;  #10 
a = 8'd170; b = 8'd77;  #10 
a = 8'd170; b = 8'd78;  #10 
a = 8'd170; b = 8'd79;  #10 
a = 8'd170; b = 8'd80;  #10 
a = 8'd170; b = 8'd81;  #10 
a = 8'd170; b = 8'd82;  #10 
a = 8'd170; b = 8'd83;  #10 
a = 8'd170; b = 8'd84;  #10 
a = 8'd170; b = 8'd85;  #10 
a = 8'd170; b = 8'd86;  #10 
a = 8'd170; b = 8'd87;  #10 
a = 8'd170; b = 8'd88;  #10 
a = 8'd170; b = 8'd89;  #10 
a = 8'd170; b = 8'd90;  #10 
a = 8'd170; b = 8'd91;  #10 
a = 8'd170; b = 8'd92;  #10 
a = 8'd170; b = 8'd93;  #10 
a = 8'd170; b = 8'd94;  #10 
a = 8'd170; b = 8'd95;  #10 
a = 8'd170; b = 8'd96;  #10 
a = 8'd170; b = 8'd97;  #10 
a = 8'd170; b = 8'd98;  #10 
a = 8'd170; b = 8'd99;  #10 
a = 8'd170; b = 8'd100;  #10 
a = 8'd170; b = 8'd101;  #10 
a = 8'd170; b = 8'd102;  #10 
a = 8'd170; b = 8'd103;  #10 
a = 8'd170; b = 8'd104;  #10 
a = 8'd170; b = 8'd105;  #10 
a = 8'd170; b = 8'd106;  #10 
a = 8'd170; b = 8'd107;  #10 
a = 8'd170; b = 8'd108;  #10 
a = 8'd170; b = 8'd109;  #10 
a = 8'd170; b = 8'd110;  #10 
a = 8'd170; b = 8'd111;  #10 
a = 8'd170; b = 8'd112;  #10 
a = 8'd170; b = 8'd113;  #10 
a = 8'd170; b = 8'd114;  #10 
a = 8'd170; b = 8'd115;  #10 
a = 8'd170; b = 8'd116;  #10 
a = 8'd170; b = 8'd117;  #10 
a = 8'd170; b = 8'd118;  #10 
a = 8'd170; b = 8'd119;  #10 
a = 8'd170; b = 8'd120;  #10 
a = 8'd170; b = 8'd121;  #10 
a = 8'd170; b = 8'd122;  #10 
a = 8'd170; b = 8'd123;  #10 
a = 8'd170; b = 8'd124;  #10 
a = 8'd170; b = 8'd125;  #10 
a = 8'd170; b = 8'd126;  #10 
a = 8'd170; b = 8'd127;  #10 
a = 8'd170; b = 8'd128;  #10 
a = 8'd170; b = 8'd129;  #10 
a = 8'd170; b = 8'd130;  #10 
a = 8'd170; b = 8'd131;  #10 
a = 8'd170; b = 8'd132;  #10 
a = 8'd170; b = 8'd133;  #10 
a = 8'd170; b = 8'd134;  #10 
a = 8'd170; b = 8'd135;  #10 
a = 8'd170; b = 8'd136;  #10 
a = 8'd170; b = 8'd137;  #10 
a = 8'd170; b = 8'd138;  #10 
a = 8'd170; b = 8'd139;  #10 
a = 8'd170; b = 8'd140;  #10 
a = 8'd170; b = 8'd141;  #10 
a = 8'd170; b = 8'd142;  #10 
a = 8'd170; b = 8'd143;  #10 
a = 8'd170; b = 8'd144;  #10 
a = 8'd170; b = 8'd145;  #10 
a = 8'd170; b = 8'd146;  #10 
a = 8'd170; b = 8'd147;  #10 
a = 8'd170; b = 8'd148;  #10 
a = 8'd170; b = 8'd149;  #10 
a = 8'd170; b = 8'd150;  #10 
a = 8'd170; b = 8'd151;  #10 
a = 8'd170; b = 8'd152;  #10 
a = 8'd170; b = 8'd153;  #10 
a = 8'd170; b = 8'd154;  #10 
a = 8'd170; b = 8'd155;  #10 
a = 8'd170; b = 8'd156;  #10 
a = 8'd170; b = 8'd157;  #10 
a = 8'd170; b = 8'd158;  #10 
a = 8'd170; b = 8'd159;  #10 
a = 8'd170; b = 8'd160;  #10 
a = 8'd170; b = 8'd161;  #10 
a = 8'd170; b = 8'd162;  #10 
a = 8'd170; b = 8'd163;  #10 
a = 8'd170; b = 8'd164;  #10 
a = 8'd170; b = 8'd165;  #10 
a = 8'd170; b = 8'd166;  #10 
a = 8'd170; b = 8'd167;  #10 
a = 8'd170; b = 8'd168;  #10 
a = 8'd170; b = 8'd169;  #10 
a = 8'd170; b = 8'd170;  #10 
a = 8'd170; b = 8'd171;  #10 
a = 8'd170; b = 8'd172;  #10 
a = 8'd170; b = 8'd173;  #10 
a = 8'd170; b = 8'd174;  #10 
a = 8'd170; b = 8'd175;  #10 
a = 8'd170; b = 8'd176;  #10 
a = 8'd170; b = 8'd177;  #10 
a = 8'd170; b = 8'd178;  #10 
a = 8'd170; b = 8'd179;  #10 
a = 8'd170; b = 8'd180;  #10 
a = 8'd170; b = 8'd181;  #10 
a = 8'd170; b = 8'd182;  #10 
a = 8'd170; b = 8'd183;  #10 
a = 8'd170; b = 8'd184;  #10 
a = 8'd170; b = 8'd185;  #10 
a = 8'd170; b = 8'd186;  #10 
a = 8'd170; b = 8'd187;  #10 
a = 8'd170; b = 8'd188;  #10 
a = 8'd170; b = 8'd189;  #10 
a = 8'd170; b = 8'd190;  #10 
a = 8'd170; b = 8'd191;  #10 
a = 8'd170; b = 8'd192;  #10 
a = 8'd170; b = 8'd193;  #10 
a = 8'd170; b = 8'd194;  #10 
a = 8'd170; b = 8'd195;  #10 
a = 8'd170; b = 8'd196;  #10 
a = 8'd170; b = 8'd197;  #10 
a = 8'd170; b = 8'd198;  #10 
a = 8'd170; b = 8'd199;  #10 
a = 8'd170; b = 8'd200;  #10 
a = 8'd170; b = 8'd201;  #10 
a = 8'd170; b = 8'd202;  #10 
a = 8'd170; b = 8'd203;  #10 
a = 8'd170; b = 8'd204;  #10 
a = 8'd170; b = 8'd205;  #10 
a = 8'd170; b = 8'd206;  #10 
a = 8'd170; b = 8'd207;  #10 
a = 8'd170; b = 8'd208;  #10 
a = 8'd170; b = 8'd209;  #10 
a = 8'd170; b = 8'd210;  #10 
a = 8'd170; b = 8'd211;  #10 
a = 8'd170; b = 8'd212;  #10 
a = 8'd170; b = 8'd213;  #10 
a = 8'd170; b = 8'd214;  #10 
a = 8'd170; b = 8'd215;  #10 
a = 8'd170; b = 8'd216;  #10 
a = 8'd170; b = 8'd217;  #10 
a = 8'd170; b = 8'd218;  #10 
a = 8'd170; b = 8'd219;  #10 
a = 8'd170; b = 8'd220;  #10 
a = 8'd170; b = 8'd221;  #10 
a = 8'd170; b = 8'd222;  #10 
a = 8'd170; b = 8'd223;  #10 
a = 8'd170; b = 8'd224;  #10 
a = 8'd170; b = 8'd225;  #10 
a = 8'd170; b = 8'd226;  #10 
a = 8'd170; b = 8'd227;  #10 
a = 8'd170; b = 8'd228;  #10 
a = 8'd170; b = 8'd229;  #10 
a = 8'd170; b = 8'd230;  #10 
a = 8'd170; b = 8'd231;  #10 
a = 8'd170; b = 8'd232;  #10 
a = 8'd170; b = 8'd233;  #10 
a = 8'd170; b = 8'd234;  #10 
a = 8'd170; b = 8'd235;  #10 
a = 8'd170; b = 8'd236;  #10 
a = 8'd170; b = 8'd237;  #10 
a = 8'd170; b = 8'd238;  #10 
a = 8'd170; b = 8'd239;  #10 
a = 8'd170; b = 8'd240;  #10 
a = 8'd170; b = 8'd241;  #10 
a = 8'd170; b = 8'd242;  #10 
a = 8'd170; b = 8'd243;  #10 
a = 8'd170; b = 8'd244;  #10 
a = 8'd170; b = 8'd245;  #10 
a = 8'd170; b = 8'd246;  #10 
a = 8'd170; b = 8'd247;  #10 
a = 8'd170; b = 8'd248;  #10 
a = 8'd170; b = 8'd249;  #10 
a = 8'd170; b = 8'd250;  #10 
a = 8'd170; b = 8'd251;  #10 
a = 8'd170; b = 8'd252;  #10 
a = 8'd170; b = 8'd253;  #10 
a = 8'd170; b = 8'd254;  #10 
a = 8'd170; b = 8'd255;  #10 
a = 8'd171; b = 8'd0;  #10 
a = 8'd171; b = 8'd1;  #10 
a = 8'd171; b = 8'd2;  #10 
a = 8'd171; b = 8'd3;  #10 
a = 8'd171; b = 8'd4;  #10 
a = 8'd171; b = 8'd5;  #10 
a = 8'd171; b = 8'd6;  #10 
a = 8'd171; b = 8'd7;  #10 
a = 8'd171; b = 8'd8;  #10 
a = 8'd171; b = 8'd9;  #10 
a = 8'd171; b = 8'd10;  #10 
a = 8'd171; b = 8'd11;  #10 
a = 8'd171; b = 8'd12;  #10 
a = 8'd171; b = 8'd13;  #10 
a = 8'd171; b = 8'd14;  #10 
a = 8'd171; b = 8'd15;  #10 
a = 8'd171; b = 8'd16;  #10 
a = 8'd171; b = 8'd17;  #10 
a = 8'd171; b = 8'd18;  #10 
a = 8'd171; b = 8'd19;  #10 
a = 8'd171; b = 8'd20;  #10 
a = 8'd171; b = 8'd21;  #10 
a = 8'd171; b = 8'd22;  #10 
a = 8'd171; b = 8'd23;  #10 
a = 8'd171; b = 8'd24;  #10 
a = 8'd171; b = 8'd25;  #10 
a = 8'd171; b = 8'd26;  #10 
a = 8'd171; b = 8'd27;  #10 
a = 8'd171; b = 8'd28;  #10 
a = 8'd171; b = 8'd29;  #10 
a = 8'd171; b = 8'd30;  #10 
a = 8'd171; b = 8'd31;  #10 
a = 8'd171; b = 8'd32;  #10 
a = 8'd171; b = 8'd33;  #10 
a = 8'd171; b = 8'd34;  #10 
a = 8'd171; b = 8'd35;  #10 
a = 8'd171; b = 8'd36;  #10 
a = 8'd171; b = 8'd37;  #10 
a = 8'd171; b = 8'd38;  #10 
a = 8'd171; b = 8'd39;  #10 
a = 8'd171; b = 8'd40;  #10 
a = 8'd171; b = 8'd41;  #10 
a = 8'd171; b = 8'd42;  #10 
a = 8'd171; b = 8'd43;  #10 
a = 8'd171; b = 8'd44;  #10 
a = 8'd171; b = 8'd45;  #10 
a = 8'd171; b = 8'd46;  #10 
a = 8'd171; b = 8'd47;  #10 
a = 8'd171; b = 8'd48;  #10 
a = 8'd171; b = 8'd49;  #10 
a = 8'd171; b = 8'd50;  #10 
a = 8'd171; b = 8'd51;  #10 
a = 8'd171; b = 8'd52;  #10 
a = 8'd171; b = 8'd53;  #10 
a = 8'd171; b = 8'd54;  #10 
a = 8'd171; b = 8'd55;  #10 
a = 8'd171; b = 8'd56;  #10 
a = 8'd171; b = 8'd57;  #10 
a = 8'd171; b = 8'd58;  #10 
a = 8'd171; b = 8'd59;  #10 
a = 8'd171; b = 8'd60;  #10 
a = 8'd171; b = 8'd61;  #10 
a = 8'd171; b = 8'd62;  #10 
a = 8'd171; b = 8'd63;  #10 
a = 8'd171; b = 8'd64;  #10 
a = 8'd171; b = 8'd65;  #10 
a = 8'd171; b = 8'd66;  #10 
a = 8'd171; b = 8'd67;  #10 
a = 8'd171; b = 8'd68;  #10 
a = 8'd171; b = 8'd69;  #10 
a = 8'd171; b = 8'd70;  #10 
a = 8'd171; b = 8'd71;  #10 
a = 8'd171; b = 8'd72;  #10 
a = 8'd171; b = 8'd73;  #10 
a = 8'd171; b = 8'd74;  #10 
a = 8'd171; b = 8'd75;  #10 
a = 8'd171; b = 8'd76;  #10 
a = 8'd171; b = 8'd77;  #10 
a = 8'd171; b = 8'd78;  #10 
a = 8'd171; b = 8'd79;  #10 
a = 8'd171; b = 8'd80;  #10 
a = 8'd171; b = 8'd81;  #10 
a = 8'd171; b = 8'd82;  #10 
a = 8'd171; b = 8'd83;  #10 
a = 8'd171; b = 8'd84;  #10 
a = 8'd171; b = 8'd85;  #10 
a = 8'd171; b = 8'd86;  #10 
a = 8'd171; b = 8'd87;  #10 
a = 8'd171; b = 8'd88;  #10 
a = 8'd171; b = 8'd89;  #10 
a = 8'd171; b = 8'd90;  #10 
a = 8'd171; b = 8'd91;  #10 
a = 8'd171; b = 8'd92;  #10 
a = 8'd171; b = 8'd93;  #10 
a = 8'd171; b = 8'd94;  #10 
a = 8'd171; b = 8'd95;  #10 
a = 8'd171; b = 8'd96;  #10 
a = 8'd171; b = 8'd97;  #10 
a = 8'd171; b = 8'd98;  #10 
a = 8'd171; b = 8'd99;  #10 
a = 8'd171; b = 8'd100;  #10 
a = 8'd171; b = 8'd101;  #10 
a = 8'd171; b = 8'd102;  #10 
a = 8'd171; b = 8'd103;  #10 
a = 8'd171; b = 8'd104;  #10 
a = 8'd171; b = 8'd105;  #10 
a = 8'd171; b = 8'd106;  #10 
a = 8'd171; b = 8'd107;  #10 
a = 8'd171; b = 8'd108;  #10 
a = 8'd171; b = 8'd109;  #10 
a = 8'd171; b = 8'd110;  #10 
a = 8'd171; b = 8'd111;  #10 
a = 8'd171; b = 8'd112;  #10 
a = 8'd171; b = 8'd113;  #10 
a = 8'd171; b = 8'd114;  #10 
a = 8'd171; b = 8'd115;  #10 
a = 8'd171; b = 8'd116;  #10 
a = 8'd171; b = 8'd117;  #10 
a = 8'd171; b = 8'd118;  #10 
a = 8'd171; b = 8'd119;  #10 
a = 8'd171; b = 8'd120;  #10 
a = 8'd171; b = 8'd121;  #10 
a = 8'd171; b = 8'd122;  #10 
a = 8'd171; b = 8'd123;  #10 
a = 8'd171; b = 8'd124;  #10 
a = 8'd171; b = 8'd125;  #10 
a = 8'd171; b = 8'd126;  #10 
a = 8'd171; b = 8'd127;  #10 
a = 8'd171; b = 8'd128;  #10 
a = 8'd171; b = 8'd129;  #10 
a = 8'd171; b = 8'd130;  #10 
a = 8'd171; b = 8'd131;  #10 
a = 8'd171; b = 8'd132;  #10 
a = 8'd171; b = 8'd133;  #10 
a = 8'd171; b = 8'd134;  #10 
a = 8'd171; b = 8'd135;  #10 
a = 8'd171; b = 8'd136;  #10 
a = 8'd171; b = 8'd137;  #10 
a = 8'd171; b = 8'd138;  #10 
a = 8'd171; b = 8'd139;  #10 
a = 8'd171; b = 8'd140;  #10 
a = 8'd171; b = 8'd141;  #10 
a = 8'd171; b = 8'd142;  #10 
a = 8'd171; b = 8'd143;  #10 
a = 8'd171; b = 8'd144;  #10 
a = 8'd171; b = 8'd145;  #10 
a = 8'd171; b = 8'd146;  #10 
a = 8'd171; b = 8'd147;  #10 
a = 8'd171; b = 8'd148;  #10 
a = 8'd171; b = 8'd149;  #10 
a = 8'd171; b = 8'd150;  #10 
a = 8'd171; b = 8'd151;  #10 
a = 8'd171; b = 8'd152;  #10 
a = 8'd171; b = 8'd153;  #10 
a = 8'd171; b = 8'd154;  #10 
a = 8'd171; b = 8'd155;  #10 
a = 8'd171; b = 8'd156;  #10 
a = 8'd171; b = 8'd157;  #10 
a = 8'd171; b = 8'd158;  #10 
a = 8'd171; b = 8'd159;  #10 
a = 8'd171; b = 8'd160;  #10 
a = 8'd171; b = 8'd161;  #10 
a = 8'd171; b = 8'd162;  #10 
a = 8'd171; b = 8'd163;  #10 
a = 8'd171; b = 8'd164;  #10 
a = 8'd171; b = 8'd165;  #10 
a = 8'd171; b = 8'd166;  #10 
a = 8'd171; b = 8'd167;  #10 
a = 8'd171; b = 8'd168;  #10 
a = 8'd171; b = 8'd169;  #10 
a = 8'd171; b = 8'd170;  #10 
a = 8'd171; b = 8'd171;  #10 
a = 8'd171; b = 8'd172;  #10 
a = 8'd171; b = 8'd173;  #10 
a = 8'd171; b = 8'd174;  #10 
a = 8'd171; b = 8'd175;  #10 
a = 8'd171; b = 8'd176;  #10 
a = 8'd171; b = 8'd177;  #10 
a = 8'd171; b = 8'd178;  #10 
a = 8'd171; b = 8'd179;  #10 
a = 8'd171; b = 8'd180;  #10 
a = 8'd171; b = 8'd181;  #10 
a = 8'd171; b = 8'd182;  #10 
a = 8'd171; b = 8'd183;  #10 
a = 8'd171; b = 8'd184;  #10 
a = 8'd171; b = 8'd185;  #10 
a = 8'd171; b = 8'd186;  #10 
a = 8'd171; b = 8'd187;  #10 
a = 8'd171; b = 8'd188;  #10 
a = 8'd171; b = 8'd189;  #10 
a = 8'd171; b = 8'd190;  #10 
a = 8'd171; b = 8'd191;  #10 
a = 8'd171; b = 8'd192;  #10 
a = 8'd171; b = 8'd193;  #10 
a = 8'd171; b = 8'd194;  #10 
a = 8'd171; b = 8'd195;  #10 
a = 8'd171; b = 8'd196;  #10 
a = 8'd171; b = 8'd197;  #10 
a = 8'd171; b = 8'd198;  #10 
a = 8'd171; b = 8'd199;  #10 
a = 8'd171; b = 8'd200;  #10 
a = 8'd171; b = 8'd201;  #10 
a = 8'd171; b = 8'd202;  #10 
a = 8'd171; b = 8'd203;  #10 
a = 8'd171; b = 8'd204;  #10 
a = 8'd171; b = 8'd205;  #10 
a = 8'd171; b = 8'd206;  #10 
a = 8'd171; b = 8'd207;  #10 
a = 8'd171; b = 8'd208;  #10 
a = 8'd171; b = 8'd209;  #10 
a = 8'd171; b = 8'd210;  #10 
a = 8'd171; b = 8'd211;  #10 
a = 8'd171; b = 8'd212;  #10 
a = 8'd171; b = 8'd213;  #10 
a = 8'd171; b = 8'd214;  #10 
a = 8'd171; b = 8'd215;  #10 
a = 8'd171; b = 8'd216;  #10 
a = 8'd171; b = 8'd217;  #10 
a = 8'd171; b = 8'd218;  #10 
a = 8'd171; b = 8'd219;  #10 
a = 8'd171; b = 8'd220;  #10 
a = 8'd171; b = 8'd221;  #10 
a = 8'd171; b = 8'd222;  #10 
a = 8'd171; b = 8'd223;  #10 
a = 8'd171; b = 8'd224;  #10 
a = 8'd171; b = 8'd225;  #10 
a = 8'd171; b = 8'd226;  #10 
a = 8'd171; b = 8'd227;  #10 
a = 8'd171; b = 8'd228;  #10 
a = 8'd171; b = 8'd229;  #10 
a = 8'd171; b = 8'd230;  #10 
a = 8'd171; b = 8'd231;  #10 
a = 8'd171; b = 8'd232;  #10 
a = 8'd171; b = 8'd233;  #10 
a = 8'd171; b = 8'd234;  #10 
a = 8'd171; b = 8'd235;  #10 
a = 8'd171; b = 8'd236;  #10 
a = 8'd171; b = 8'd237;  #10 
a = 8'd171; b = 8'd238;  #10 
a = 8'd171; b = 8'd239;  #10 
a = 8'd171; b = 8'd240;  #10 
a = 8'd171; b = 8'd241;  #10 
a = 8'd171; b = 8'd242;  #10 
a = 8'd171; b = 8'd243;  #10 
a = 8'd171; b = 8'd244;  #10 
a = 8'd171; b = 8'd245;  #10 
a = 8'd171; b = 8'd246;  #10 
a = 8'd171; b = 8'd247;  #10 
a = 8'd171; b = 8'd248;  #10 
a = 8'd171; b = 8'd249;  #10 
a = 8'd171; b = 8'd250;  #10 
a = 8'd171; b = 8'd251;  #10 
a = 8'd171; b = 8'd252;  #10 
a = 8'd171; b = 8'd253;  #10 
a = 8'd171; b = 8'd254;  #10 
a = 8'd171; b = 8'd255;  #10 
a = 8'd172; b = 8'd0;  #10 
a = 8'd172; b = 8'd1;  #10 
a = 8'd172; b = 8'd2;  #10 
a = 8'd172; b = 8'd3;  #10 
a = 8'd172; b = 8'd4;  #10 
a = 8'd172; b = 8'd5;  #10 
a = 8'd172; b = 8'd6;  #10 
a = 8'd172; b = 8'd7;  #10 
a = 8'd172; b = 8'd8;  #10 
a = 8'd172; b = 8'd9;  #10 
a = 8'd172; b = 8'd10;  #10 
a = 8'd172; b = 8'd11;  #10 
a = 8'd172; b = 8'd12;  #10 
a = 8'd172; b = 8'd13;  #10 
a = 8'd172; b = 8'd14;  #10 
a = 8'd172; b = 8'd15;  #10 
a = 8'd172; b = 8'd16;  #10 
a = 8'd172; b = 8'd17;  #10 
a = 8'd172; b = 8'd18;  #10 
a = 8'd172; b = 8'd19;  #10 
a = 8'd172; b = 8'd20;  #10 
a = 8'd172; b = 8'd21;  #10 
a = 8'd172; b = 8'd22;  #10 
a = 8'd172; b = 8'd23;  #10 
a = 8'd172; b = 8'd24;  #10 
a = 8'd172; b = 8'd25;  #10 
a = 8'd172; b = 8'd26;  #10 
a = 8'd172; b = 8'd27;  #10 
a = 8'd172; b = 8'd28;  #10 
a = 8'd172; b = 8'd29;  #10 
a = 8'd172; b = 8'd30;  #10 
a = 8'd172; b = 8'd31;  #10 
a = 8'd172; b = 8'd32;  #10 
a = 8'd172; b = 8'd33;  #10 
a = 8'd172; b = 8'd34;  #10 
a = 8'd172; b = 8'd35;  #10 
a = 8'd172; b = 8'd36;  #10 
a = 8'd172; b = 8'd37;  #10 
a = 8'd172; b = 8'd38;  #10 
a = 8'd172; b = 8'd39;  #10 
a = 8'd172; b = 8'd40;  #10 
a = 8'd172; b = 8'd41;  #10 
a = 8'd172; b = 8'd42;  #10 
a = 8'd172; b = 8'd43;  #10 
a = 8'd172; b = 8'd44;  #10 
a = 8'd172; b = 8'd45;  #10 
a = 8'd172; b = 8'd46;  #10 
a = 8'd172; b = 8'd47;  #10 
a = 8'd172; b = 8'd48;  #10 
a = 8'd172; b = 8'd49;  #10 
a = 8'd172; b = 8'd50;  #10 
a = 8'd172; b = 8'd51;  #10 
a = 8'd172; b = 8'd52;  #10 
a = 8'd172; b = 8'd53;  #10 
a = 8'd172; b = 8'd54;  #10 
a = 8'd172; b = 8'd55;  #10 
a = 8'd172; b = 8'd56;  #10 
a = 8'd172; b = 8'd57;  #10 
a = 8'd172; b = 8'd58;  #10 
a = 8'd172; b = 8'd59;  #10 
a = 8'd172; b = 8'd60;  #10 
a = 8'd172; b = 8'd61;  #10 
a = 8'd172; b = 8'd62;  #10 
a = 8'd172; b = 8'd63;  #10 
a = 8'd172; b = 8'd64;  #10 
a = 8'd172; b = 8'd65;  #10 
a = 8'd172; b = 8'd66;  #10 
a = 8'd172; b = 8'd67;  #10 
a = 8'd172; b = 8'd68;  #10 
a = 8'd172; b = 8'd69;  #10 
a = 8'd172; b = 8'd70;  #10 
a = 8'd172; b = 8'd71;  #10 
a = 8'd172; b = 8'd72;  #10 
a = 8'd172; b = 8'd73;  #10 
a = 8'd172; b = 8'd74;  #10 
a = 8'd172; b = 8'd75;  #10 
a = 8'd172; b = 8'd76;  #10 
a = 8'd172; b = 8'd77;  #10 
a = 8'd172; b = 8'd78;  #10 
a = 8'd172; b = 8'd79;  #10 
a = 8'd172; b = 8'd80;  #10 
a = 8'd172; b = 8'd81;  #10 
a = 8'd172; b = 8'd82;  #10 
a = 8'd172; b = 8'd83;  #10 
a = 8'd172; b = 8'd84;  #10 
a = 8'd172; b = 8'd85;  #10 
a = 8'd172; b = 8'd86;  #10 
a = 8'd172; b = 8'd87;  #10 
a = 8'd172; b = 8'd88;  #10 
a = 8'd172; b = 8'd89;  #10 
a = 8'd172; b = 8'd90;  #10 
a = 8'd172; b = 8'd91;  #10 
a = 8'd172; b = 8'd92;  #10 
a = 8'd172; b = 8'd93;  #10 
a = 8'd172; b = 8'd94;  #10 
a = 8'd172; b = 8'd95;  #10 
a = 8'd172; b = 8'd96;  #10 
a = 8'd172; b = 8'd97;  #10 
a = 8'd172; b = 8'd98;  #10 
a = 8'd172; b = 8'd99;  #10 
a = 8'd172; b = 8'd100;  #10 
a = 8'd172; b = 8'd101;  #10 
a = 8'd172; b = 8'd102;  #10 
a = 8'd172; b = 8'd103;  #10 
a = 8'd172; b = 8'd104;  #10 
a = 8'd172; b = 8'd105;  #10 
a = 8'd172; b = 8'd106;  #10 
a = 8'd172; b = 8'd107;  #10 
a = 8'd172; b = 8'd108;  #10 
a = 8'd172; b = 8'd109;  #10 
a = 8'd172; b = 8'd110;  #10 
a = 8'd172; b = 8'd111;  #10 
a = 8'd172; b = 8'd112;  #10 
a = 8'd172; b = 8'd113;  #10 
a = 8'd172; b = 8'd114;  #10 
a = 8'd172; b = 8'd115;  #10 
a = 8'd172; b = 8'd116;  #10 
a = 8'd172; b = 8'd117;  #10 
a = 8'd172; b = 8'd118;  #10 
a = 8'd172; b = 8'd119;  #10 
a = 8'd172; b = 8'd120;  #10 
a = 8'd172; b = 8'd121;  #10 
a = 8'd172; b = 8'd122;  #10 
a = 8'd172; b = 8'd123;  #10 
a = 8'd172; b = 8'd124;  #10 
a = 8'd172; b = 8'd125;  #10 
a = 8'd172; b = 8'd126;  #10 
a = 8'd172; b = 8'd127;  #10 
a = 8'd172; b = 8'd128;  #10 
a = 8'd172; b = 8'd129;  #10 
a = 8'd172; b = 8'd130;  #10 
a = 8'd172; b = 8'd131;  #10 
a = 8'd172; b = 8'd132;  #10 
a = 8'd172; b = 8'd133;  #10 
a = 8'd172; b = 8'd134;  #10 
a = 8'd172; b = 8'd135;  #10 
a = 8'd172; b = 8'd136;  #10 
a = 8'd172; b = 8'd137;  #10 
a = 8'd172; b = 8'd138;  #10 
a = 8'd172; b = 8'd139;  #10 
a = 8'd172; b = 8'd140;  #10 
a = 8'd172; b = 8'd141;  #10 
a = 8'd172; b = 8'd142;  #10 
a = 8'd172; b = 8'd143;  #10 
a = 8'd172; b = 8'd144;  #10 
a = 8'd172; b = 8'd145;  #10 
a = 8'd172; b = 8'd146;  #10 
a = 8'd172; b = 8'd147;  #10 
a = 8'd172; b = 8'd148;  #10 
a = 8'd172; b = 8'd149;  #10 
a = 8'd172; b = 8'd150;  #10 
a = 8'd172; b = 8'd151;  #10 
a = 8'd172; b = 8'd152;  #10 
a = 8'd172; b = 8'd153;  #10 
a = 8'd172; b = 8'd154;  #10 
a = 8'd172; b = 8'd155;  #10 
a = 8'd172; b = 8'd156;  #10 
a = 8'd172; b = 8'd157;  #10 
a = 8'd172; b = 8'd158;  #10 
a = 8'd172; b = 8'd159;  #10 
a = 8'd172; b = 8'd160;  #10 
a = 8'd172; b = 8'd161;  #10 
a = 8'd172; b = 8'd162;  #10 
a = 8'd172; b = 8'd163;  #10 
a = 8'd172; b = 8'd164;  #10 
a = 8'd172; b = 8'd165;  #10 
a = 8'd172; b = 8'd166;  #10 
a = 8'd172; b = 8'd167;  #10 
a = 8'd172; b = 8'd168;  #10 
a = 8'd172; b = 8'd169;  #10 
a = 8'd172; b = 8'd170;  #10 
a = 8'd172; b = 8'd171;  #10 
a = 8'd172; b = 8'd172;  #10 
a = 8'd172; b = 8'd173;  #10 
a = 8'd172; b = 8'd174;  #10 
a = 8'd172; b = 8'd175;  #10 
a = 8'd172; b = 8'd176;  #10 
a = 8'd172; b = 8'd177;  #10 
a = 8'd172; b = 8'd178;  #10 
a = 8'd172; b = 8'd179;  #10 
a = 8'd172; b = 8'd180;  #10 
a = 8'd172; b = 8'd181;  #10 
a = 8'd172; b = 8'd182;  #10 
a = 8'd172; b = 8'd183;  #10 
a = 8'd172; b = 8'd184;  #10 
a = 8'd172; b = 8'd185;  #10 
a = 8'd172; b = 8'd186;  #10 
a = 8'd172; b = 8'd187;  #10 
a = 8'd172; b = 8'd188;  #10 
a = 8'd172; b = 8'd189;  #10 
a = 8'd172; b = 8'd190;  #10 
a = 8'd172; b = 8'd191;  #10 
a = 8'd172; b = 8'd192;  #10 
a = 8'd172; b = 8'd193;  #10 
a = 8'd172; b = 8'd194;  #10 
a = 8'd172; b = 8'd195;  #10 
a = 8'd172; b = 8'd196;  #10 
a = 8'd172; b = 8'd197;  #10 
a = 8'd172; b = 8'd198;  #10 
a = 8'd172; b = 8'd199;  #10 
a = 8'd172; b = 8'd200;  #10 
a = 8'd172; b = 8'd201;  #10 
a = 8'd172; b = 8'd202;  #10 
a = 8'd172; b = 8'd203;  #10 
a = 8'd172; b = 8'd204;  #10 
a = 8'd172; b = 8'd205;  #10 
a = 8'd172; b = 8'd206;  #10 
a = 8'd172; b = 8'd207;  #10 
a = 8'd172; b = 8'd208;  #10 
a = 8'd172; b = 8'd209;  #10 
a = 8'd172; b = 8'd210;  #10 
a = 8'd172; b = 8'd211;  #10 
a = 8'd172; b = 8'd212;  #10 
a = 8'd172; b = 8'd213;  #10 
a = 8'd172; b = 8'd214;  #10 
a = 8'd172; b = 8'd215;  #10 
a = 8'd172; b = 8'd216;  #10 
a = 8'd172; b = 8'd217;  #10 
a = 8'd172; b = 8'd218;  #10 
a = 8'd172; b = 8'd219;  #10 
a = 8'd172; b = 8'd220;  #10 
a = 8'd172; b = 8'd221;  #10 
a = 8'd172; b = 8'd222;  #10 
a = 8'd172; b = 8'd223;  #10 
a = 8'd172; b = 8'd224;  #10 
a = 8'd172; b = 8'd225;  #10 
a = 8'd172; b = 8'd226;  #10 
a = 8'd172; b = 8'd227;  #10 
a = 8'd172; b = 8'd228;  #10 
a = 8'd172; b = 8'd229;  #10 
a = 8'd172; b = 8'd230;  #10 
a = 8'd172; b = 8'd231;  #10 
a = 8'd172; b = 8'd232;  #10 
a = 8'd172; b = 8'd233;  #10 
a = 8'd172; b = 8'd234;  #10 
a = 8'd172; b = 8'd235;  #10 
a = 8'd172; b = 8'd236;  #10 
a = 8'd172; b = 8'd237;  #10 
a = 8'd172; b = 8'd238;  #10 
a = 8'd172; b = 8'd239;  #10 
a = 8'd172; b = 8'd240;  #10 
a = 8'd172; b = 8'd241;  #10 
a = 8'd172; b = 8'd242;  #10 
a = 8'd172; b = 8'd243;  #10 
a = 8'd172; b = 8'd244;  #10 
a = 8'd172; b = 8'd245;  #10 
a = 8'd172; b = 8'd246;  #10 
a = 8'd172; b = 8'd247;  #10 
a = 8'd172; b = 8'd248;  #10 
a = 8'd172; b = 8'd249;  #10 
a = 8'd172; b = 8'd250;  #10 
a = 8'd172; b = 8'd251;  #10 
a = 8'd172; b = 8'd252;  #10 
a = 8'd172; b = 8'd253;  #10 
a = 8'd172; b = 8'd254;  #10 
a = 8'd172; b = 8'd255;  #10 
a = 8'd173; b = 8'd0;  #10 
a = 8'd173; b = 8'd1;  #10 
a = 8'd173; b = 8'd2;  #10 
a = 8'd173; b = 8'd3;  #10 
a = 8'd173; b = 8'd4;  #10 
a = 8'd173; b = 8'd5;  #10 
a = 8'd173; b = 8'd6;  #10 
a = 8'd173; b = 8'd7;  #10 
a = 8'd173; b = 8'd8;  #10 
a = 8'd173; b = 8'd9;  #10 
a = 8'd173; b = 8'd10;  #10 
a = 8'd173; b = 8'd11;  #10 
a = 8'd173; b = 8'd12;  #10 
a = 8'd173; b = 8'd13;  #10 
a = 8'd173; b = 8'd14;  #10 
a = 8'd173; b = 8'd15;  #10 
a = 8'd173; b = 8'd16;  #10 
a = 8'd173; b = 8'd17;  #10 
a = 8'd173; b = 8'd18;  #10 
a = 8'd173; b = 8'd19;  #10 
a = 8'd173; b = 8'd20;  #10 
a = 8'd173; b = 8'd21;  #10 
a = 8'd173; b = 8'd22;  #10 
a = 8'd173; b = 8'd23;  #10 
a = 8'd173; b = 8'd24;  #10 
a = 8'd173; b = 8'd25;  #10 
a = 8'd173; b = 8'd26;  #10 
a = 8'd173; b = 8'd27;  #10 
a = 8'd173; b = 8'd28;  #10 
a = 8'd173; b = 8'd29;  #10 
a = 8'd173; b = 8'd30;  #10 
a = 8'd173; b = 8'd31;  #10 
a = 8'd173; b = 8'd32;  #10 
a = 8'd173; b = 8'd33;  #10 
a = 8'd173; b = 8'd34;  #10 
a = 8'd173; b = 8'd35;  #10 
a = 8'd173; b = 8'd36;  #10 
a = 8'd173; b = 8'd37;  #10 
a = 8'd173; b = 8'd38;  #10 
a = 8'd173; b = 8'd39;  #10 
a = 8'd173; b = 8'd40;  #10 
a = 8'd173; b = 8'd41;  #10 
a = 8'd173; b = 8'd42;  #10 
a = 8'd173; b = 8'd43;  #10 
a = 8'd173; b = 8'd44;  #10 
a = 8'd173; b = 8'd45;  #10 
a = 8'd173; b = 8'd46;  #10 
a = 8'd173; b = 8'd47;  #10 
a = 8'd173; b = 8'd48;  #10 
a = 8'd173; b = 8'd49;  #10 
a = 8'd173; b = 8'd50;  #10 
a = 8'd173; b = 8'd51;  #10 
a = 8'd173; b = 8'd52;  #10 
a = 8'd173; b = 8'd53;  #10 
a = 8'd173; b = 8'd54;  #10 
a = 8'd173; b = 8'd55;  #10 
a = 8'd173; b = 8'd56;  #10 
a = 8'd173; b = 8'd57;  #10 
a = 8'd173; b = 8'd58;  #10 
a = 8'd173; b = 8'd59;  #10 
a = 8'd173; b = 8'd60;  #10 
a = 8'd173; b = 8'd61;  #10 
a = 8'd173; b = 8'd62;  #10 
a = 8'd173; b = 8'd63;  #10 
a = 8'd173; b = 8'd64;  #10 
a = 8'd173; b = 8'd65;  #10 
a = 8'd173; b = 8'd66;  #10 
a = 8'd173; b = 8'd67;  #10 
a = 8'd173; b = 8'd68;  #10 
a = 8'd173; b = 8'd69;  #10 
a = 8'd173; b = 8'd70;  #10 
a = 8'd173; b = 8'd71;  #10 
a = 8'd173; b = 8'd72;  #10 
a = 8'd173; b = 8'd73;  #10 
a = 8'd173; b = 8'd74;  #10 
a = 8'd173; b = 8'd75;  #10 
a = 8'd173; b = 8'd76;  #10 
a = 8'd173; b = 8'd77;  #10 
a = 8'd173; b = 8'd78;  #10 
a = 8'd173; b = 8'd79;  #10 
a = 8'd173; b = 8'd80;  #10 
a = 8'd173; b = 8'd81;  #10 
a = 8'd173; b = 8'd82;  #10 
a = 8'd173; b = 8'd83;  #10 
a = 8'd173; b = 8'd84;  #10 
a = 8'd173; b = 8'd85;  #10 
a = 8'd173; b = 8'd86;  #10 
a = 8'd173; b = 8'd87;  #10 
a = 8'd173; b = 8'd88;  #10 
a = 8'd173; b = 8'd89;  #10 
a = 8'd173; b = 8'd90;  #10 
a = 8'd173; b = 8'd91;  #10 
a = 8'd173; b = 8'd92;  #10 
a = 8'd173; b = 8'd93;  #10 
a = 8'd173; b = 8'd94;  #10 
a = 8'd173; b = 8'd95;  #10 
a = 8'd173; b = 8'd96;  #10 
a = 8'd173; b = 8'd97;  #10 
a = 8'd173; b = 8'd98;  #10 
a = 8'd173; b = 8'd99;  #10 
a = 8'd173; b = 8'd100;  #10 
a = 8'd173; b = 8'd101;  #10 
a = 8'd173; b = 8'd102;  #10 
a = 8'd173; b = 8'd103;  #10 
a = 8'd173; b = 8'd104;  #10 
a = 8'd173; b = 8'd105;  #10 
a = 8'd173; b = 8'd106;  #10 
a = 8'd173; b = 8'd107;  #10 
a = 8'd173; b = 8'd108;  #10 
a = 8'd173; b = 8'd109;  #10 
a = 8'd173; b = 8'd110;  #10 
a = 8'd173; b = 8'd111;  #10 
a = 8'd173; b = 8'd112;  #10 
a = 8'd173; b = 8'd113;  #10 
a = 8'd173; b = 8'd114;  #10 
a = 8'd173; b = 8'd115;  #10 
a = 8'd173; b = 8'd116;  #10 
a = 8'd173; b = 8'd117;  #10 
a = 8'd173; b = 8'd118;  #10 
a = 8'd173; b = 8'd119;  #10 
a = 8'd173; b = 8'd120;  #10 
a = 8'd173; b = 8'd121;  #10 
a = 8'd173; b = 8'd122;  #10 
a = 8'd173; b = 8'd123;  #10 
a = 8'd173; b = 8'd124;  #10 
a = 8'd173; b = 8'd125;  #10 
a = 8'd173; b = 8'd126;  #10 
a = 8'd173; b = 8'd127;  #10 
a = 8'd173; b = 8'd128;  #10 
a = 8'd173; b = 8'd129;  #10 
a = 8'd173; b = 8'd130;  #10 
a = 8'd173; b = 8'd131;  #10 
a = 8'd173; b = 8'd132;  #10 
a = 8'd173; b = 8'd133;  #10 
a = 8'd173; b = 8'd134;  #10 
a = 8'd173; b = 8'd135;  #10 
a = 8'd173; b = 8'd136;  #10 
a = 8'd173; b = 8'd137;  #10 
a = 8'd173; b = 8'd138;  #10 
a = 8'd173; b = 8'd139;  #10 
a = 8'd173; b = 8'd140;  #10 
a = 8'd173; b = 8'd141;  #10 
a = 8'd173; b = 8'd142;  #10 
a = 8'd173; b = 8'd143;  #10 
a = 8'd173; b = 8'd144;  #10 
a = 8'd173; b = 8'd145;  #10 
a = 8'd173; b = 8'd146;  #10 
a = 8'd173; b = 8'd147;  #10 
a = 8'd173; b = 8'd148;  #10 
a = 8'd173; b = 8'd149;  #10 
a = 8'd173; b = 8'd150;  #10 
a = 8'd173; b = 8'd151;  #10 
a = 8'd173; b = 8'd152;  #10 
a = 8'd173; b = 8'd153;  #10 
a = 8'd173; b = 8'd154;  #10 
a = 8'd173; b = 8'd155;  #10 
a = 8'd173; b = 8'd156;  #10 
a = 8'd173; b = 8'd157;  #10 
a = 8'd173; b = 8'd158;  #10 
a = 8'd173; b = 8'd159;  #10 
a = 8'd173; b = 8'd160;  #10 
a = 8'd173; b = 8'd161;  #10 
a = 8'd173; b = 8'd162;  #10 
a = 8'd173; b = 8'd163;  #10 
a = 8'd173; b = 8'd164;  #10 
a = 8'd173; b = 8'd165;  #10 
a = 8'd173; b = 8'd166;  #10 
a = 8'd173; b = 8'd167;  #10 
a = 8'd173; b = 8'd168;  #10 
a = 8'd173; b = 8'd169;  #10 
a = 8'd173; b = 8'd170;  #10 
a = 8'd173; b = 8'd171;  #10 
a = 8'd173; b = 8'd172;  #10 
a = 8'd173; b = 8'd173;  #10 
a = 8'd173; b = 8'd174;  #10 
a = 8'd173; b = 8'd175;  #10 
a = 8'd173; b = 8'd176;  #10 
a = 8'd173; b = 8'd177;  #10 
a = 8'd173; b = 8'd178;  #10 
a = 8'd173; b = 8'd179;  #10 
a = 8'd173; b = 8'd180;  #10 
a = 8'd173; b = 8'd181;  #10 
a = 8'd173; b = 8'd182;  #10 
a = 8'd173; b = 8'd183;  #10 
a = 8'd173; b = 8'd184;  #10 
a = 8'd173; b = 8'd185;  #10 
a = 8'd173; b = 8'd186;  #10 
a = 8'd173; b = 8'd187;  #10 
a = 8'd173; b = 8'd188;  #10 
a = 8'd173; b = 8'd189;  #10 
a = 8'd173; b = 8'd190;  #10 
a = 8'd173; b = 8'd191;  #10 
a = 8'd173; b = 8'd192;  #10 
a = 8'd173; b = 8'd193;  #10 
a = 8'd173; b = 8'd194;  #10 
a = 8'd173; b = 8'd195;  #10 
a = 8'd173; b = 8'd196;  #10 
a = 8'd173; b = 8'd197;  #10 
a = 8'd173; b = 8'd198;  #10 
a = 8'd173; b = 8'd199;  #10 
a = 8'd173; b = 8'd200;  #10 
a = 8'd173; b = 8'd201;  #10 
a = 8'd173; b = 8'd202;  #10 
a = 8'd173; b = 8'd203;  #10 
a = 8'd173; b = 8'd204;  #10 
a = 8'd173; b = 8'd205;  #10 
a = 8'd173; b = 8'd206;  #10 
a = 8'd173; b = 8'd207;  #10 
a = 8'd173; b = 8'd208;  #10 
a = 8'd173; b = 8'd209;  #10 
a = 8'd173; b = 8'd210;  #10 
a = 8'd173; b = 8'd211;  #10 
a = 8'd173; b = 8'd212;  #10 
a = 8'd173; b = 8'd213;  #10 
a = 8'd173; b = 8'd214;  #10 
a = 8'd173; b = 8'd215;  #10 
a = 8'd173; b = 8'd216;  #10 
a = 8'd173; b = 8'd217;  #10 
a = 8'd173; b = 8'd218;  #10 
a = 8'd173; b = 8'd219;  #10 
a = 8'd173; b = 8'd220;  #10 
a = 8'd173; b = 8'd221;  #10 
a = 8'd173; b = 8'd222;  #10 
a = 8'd173; b = 8'd223;  #10 
a = 8'd173; b = 8'd224;  #10 
a = 8'd173; b = 8'd225;  #10 
a = 8'd173; b = 8'd226;  #10 
a = 8'd173; b = 8'd227;  #10 
a = 8'd173; b = 8'd228;  #10 
a = 8'd173; b = 8'd229;  #10 
a = 8'd173; b = 8'd230;  #10 
a = 8'd173; b = 8'd231;  #10 
a = 8'd173; b = 8'd232;  #10 
a = 8'd173; b = 8'd233;  #10 
a = 8'd173; b = 8'd234;  #10 
a = 8'd173; b = 8'd235;  #10 
a = 8'd173; b = 8'd236;  #10 
a = 8'd173; b = 8'd237;  #10 
a = 8'd173; b = 8'd238;  #10 
a = 8'd173; b = 8'd239;  #10 
a = 8'd173; b = 8'd240;  #10 
a = 8'd173; b = 8'd241;  #10 
a = 8'd173; b = 8'd242;  #10 
a = 8'd173; b = 8'd243;  #10 
a = 8'd173; b = 8'd244;  #10 
a = 8'd173; b = 8'd245;  #10 
a = 8'd173; b = 8'd246;  #10 
a = 8'd173; b = 8'd247;  #10 
a = 8'd173; b = 8'd248;  #10 
a = 8'd173; b = 8'd249;  #10 
a = 8'd173; b = 8'd250;  #10 
a = 8'd173; b = 8'd251;  #10 
a = 8'd173; b = 8'd252;  #10 
a = 8'd173; b = 8'd253;  #10 
a = 8'd173; b = 8'd254;  #10 
a = 8'd173; b = 8'd255;  #10 
a = 8'd174; b = 8'd0;  #10 
a = 8'd174; b = 8'd1;  #10 
a = 8'd174; b = 8'd2;  #10 
a = 8'd174; b = 8'd3;  #10 
a = 8'd174; b = 8'd4;  #10 
a = 8'd174; b = 8'd5;  #10 
a = 8'd174; b = 8'd6;  #10 
a = 8'd174; b = 8'd7;  #10 
a = 8'd174; b = 8'd8;  #10 
a = 8'd174; b = 8'd9;  #10 
a = 8'd174; b = 8'd10;  #10 
a = 8'd174; b = 8'd11;  #10 
a = 8'd174; b = 8'd12;  #10 
a = 8'd174; b = 8'd13;  #10 
a = 8'd174; b = 8'd14;  #10 
a = 8'd174; b = 8'd15;  #10 
a = 8'd174; b = 8'd16;  #10 
a = 8'd174; b = 8'd17;  #10 
a = 8'd174; b = 8'd18;  #10 
a = 8'd174; b = 8'd19;  #10 
a = 8'd174; b = 8'd20;  #10 
a = 8'd174; b = 8'd21;  #10 
a = 8'd174; b = 8'd22;  #10 
a = 8'd174; b = 8'd23;  #10 
a = 8'd174; b = 8'd24;  #10 
a = 8'd174; b = 8'd25;  #10 
a = 8'd174; b = 8'd26;  #10 
a = 8'd174; b = 8'd27;  #10 
a = 8'd174; b = 8'd28;  #10 
a = 8'd174; b = 8'd29;  #10 
a = 8'd174; b = 8'd30;  #10 
a = 8'd174; b = 8'd31;  #10 
a = 8'd174; b = 8'd32;  #10 
a = 8'd174; b = 8'd33;  #10 
a = 8'd174; b = 8'd34;  #10 
a = 8'd174; b = 8'd35;  #10 
a = 8'd174; b = 8'd36;  #10 
a = 8'd174; b = 8'd37;  #10 
a = 8'd174; b = 8'd38;  #10 
a = 8'd174; b = 8'd39;  #10 
a = 8'd174; b = 8'd40;  #10 
a = 8'd174; b = 8'd41;  #10 
a = 8'd174; b = 8'd42;  #10 
a = 8'd174; b = 8'd43;  #10 
a = 8'd174; b = 8'd44;  #10 
a = 8'd174; b = 8'd45;  #10 
a = 8'd174; b = 8'd46;  #10 
a = 8'd174; b = 8'd47;  #10 
a = 8'd174; b = 8'd48;  #10 
a = 8'd174; b = 8'd49;  #10 
a = 8'd174; b = 8'd50;  #10 
a = 8'd174; b = 8'd51;  #10 
a = 8'd174; b = 8'd52;  #10 
a = 8'd174; b = 8'd53;  #10 
a = 8'd174; b = 8'd54;  #10 
a = 8'd174; b = 8'd55;  #10 
a = 8'd174; b = 8'd56;  #10 
a = 8'd174; b = 8'd57;  #10 
a = 8'd174; b = 8'd58;  #10 
a = 8'd174; b = 8'd59;  #10 
a = 8'd174; b = 8'd60;  #10 
a = 8'd174; b = 8'd61;  #10 
a = 8'd174; b = 8'd62;  #10 
a = 8'd174; b = 8'd63;  #10 
a = 8'd174; b = 8'd64;  #10 
a = 8'd174; b = 8'd65;  #10 
a = 8'd174; b = 8'd66;  #10 
a = 8'd174; b = 8'd67;  #10 
a = 8'd174; b = 8'd68;  #10 
a = 8'd174; b = 8'd69;  #10 
a = 8'd174; b = 8'd70;  #10 
a = 8'd174; b = 8'd71;  #10 
a = 8'd174; b = 8'd72;  #10 
a = 8'd174; b = 8'd73;  #10 
a = 8'd174; b = 8'd74;  #10 
a = 8'd174; b = 8'd75;  #10 
a = 8'd174; b = 8'd76;  #10 
a = 8'd174; b = 8'd77;  #10 
a = 8'd174; b = 8'd78;  #10 
a = 8'd174; b = 8'd79;  #10 
a = 8'd174; b = 8'd80;  #10 
a = 8'd174; b = 8'd81;  #10 
a = 8'd174; b = 8'd82;  #10 
a = 8'd174; b = 8'd83;  #10 
a = 8'd174; b = 8'd84;  #10 
a = 8'd174; b = 8'd85;  #10 
a = 8'd174; b = 8'd86;  #10 
a = 8'd174; b = 8'd87;  #10 
a = 8'd174; b = 8'd88;  #10 
a = 8'd174; b = 8'd89;  #10 
a = 8'd174; b = 8'd90;  #10 
a = 8'd174; b = 8'd91;  #10 
a = 8'd174; b = 8'd92;  #10 
a = 8'd174; b = 8'd93;  #10 
a = 8'd174; b = 8'd94;  #10 
a = 8'd174; b = 8'd95;  #10 
a = 8'd174; b = 8'd96;  #10 
a = 8'd174; b = 8'd97;  #10 
a = 8'd174; b = 8'd98;  #10 
a = 8'd174; b = 8'd99;  #10 
a = 8'd174; b = 8'd100;  #10 
a = 8'd174; b = 8'd101;  #10 
a = 8'd174; b = 8'd102;  #10 
a = 8'd174; b = 8'd103;  #10 
a = 8'd174; b = 8'd104;  #10 
a = 8'd174; b = 8'd105;  #10 
a = 8'd174; b = 8'd106;  #10 
a = 8'd174; b = 8'd107;  #10 
a = 8'd174; b = 8'd108;  #10 
a = 8'd174; b = 8'd109;  #10 
a = 8'd174; b = 8'd110;  #10 
a = 8'd174; b = 8'd111;  #10 
a = 8'd174; b = 8'd112;  #10 
a = 8'd174; b = 8'd113;  #10 
a = 8'd174; b = 8'd114;  #10 
a = 8'd174; b = 8'd115;  #10 
a = 8'd174; b = 8'd116;  #10 
a = 8'd174; b = 8'd117;  #10 
a = 8'd174; b = 8'd118;  #10 
a = 8'd174; b = 8'd119;  #10 
a = 8'd174; b = 8'd120;  #10 
a = 8'd174; b = 8'd121;  #10 
a = 8'd174; b = 8'd122;  #10 
a = 8'd174; b = 8'd123;  #10 
a = 8'd174; b = 8'd124;  #10 
a = 8'd174; b = 8'd125;  #10 
a = 8'd174; b = 8'd126;  #10 
a = 8'd174; b = 8'd127;  #10 
a = 8'd174; b = 8'd128;  #10 
a = 8'd174; b = 8'd129;  #10 
a = 8'd174; b = 8'd130;  #10 
a = 8'd174; b = 8'd131;  #10 
a = 8'd174; b = 8'd132;  #10 
a = 8'd174; b = 8'd133;  #10 
a = 8'd174; b = 8'd134;  #10 
a = 8'd174; b = 8'd135;  #10 
a = 8'd174; b = 8'd136;  #10 
a = 8'd174; b = 8'd137;  #10 
a = 8'd174; b = 8'd138;  #10 
a = 8'd174; b = 8'd139;  #10 
a = 8'd174; b = 8'd140;  #10 
a = 8'd174; b = 8'd141;  #10 
a = 8'd174; b = 8'd142;  #10 
a = 8'd174; b = 8'd143;  #10 
a = 8'd174; b = 8'd144;  #10 
a = 8'd174; b = 8'd145;  #10 
a = 8'd174; b = 8'd146;  #10 
a = 8'd174; b = 8'd147;  #10 
a = 8'd174; b = 8'd148;  #10 
a = 8'd174; b = 8'd149;  #10 
a = 8'd174; b = 8'd150;  #10 
a = 8'd174; b = 8'd151;  #10 
a = 8'd174; b = 8'd152;  #10 
a = 8'd174; b = 8'd153;  #10 
a = 8'd174; b = 8'd154;  #10 
a = 8'd174; b = 8'd155;  #10 
a = 8'd174; b = 8'd156;  #10 
a = 8'd174; b = 8'd157;  #10 
a = 8'd174; b = 8'd158;  #10 
a = 8'd174; b = 8'd159;  #10 
a = 8'd174; b = 8'd160;  #10 
a = 8'd174; b = 8'd161;  #10 
a = 8'd174; b = 8'd162;  #10 
a = 8'd174; b = 8'd163;  #10 
a = 8'd174; b = 8'd164;  #10 
a = 8'd174; b = 8'd165;  #10 
a = 8'd174; b = 8'd166;  #10 
a = 8'd174; b = 8'd167;  #10 
a = 8'd174; b = 8'd168;  #10 
a = 8'd174; b = 8'd169;  #10 
a = 8'd174; b = 8'd170;  #10 
a = 8'd174; b = 8'd171;  #10 
a = 8'd174; b = 8'd172;  #10 
a = 8'd174; b = 8'd173;  #10 
a = 8'd174; b = 8'd174;  #10 
a = 8'd174; b = 8'd175;  #10 
a = 8'd174; b = 8'd176;  #10 
a = 8'd174; b = 8'd177;  #10 
a = 8'd174; b = 8'd178;  #10 
a = 8'd174; b = 8'd179;  #10 
a = 8'd174; b = 8'd180;  #10 
a = 8'd174; b = 8'd181;  #10 
a = 8'd174; b = 8'd182;  #10 
a = 8'd174; b = 8'd183;  #10 
a = 8'd174; b = 8'd184;  #10 
a = 8'd174; b = 8'd185;  #10 
a = 8'd174; b = 8'd186;  #10 
a = 8'd174; b = 8'd187;  #10 
a = 8'd174; b = 8'd188;  #10 
a = 8'd174; b = 8'd189;  #10 
a = 8'd174; b = 8'd190;  #10 
a = 8'd174; b = 8'd191;  #10 
a = 8'd174; b = 8'd192;  #10 
a = 8'd174; b = 8'd193;  #10 
a = 8'd174; b = 8'd194;  #10 
a = 8'd174; b = 8'd195;  #10 
a = 8'd174; b = 8'd196;  #10 
a = 8'd174; b = 8'd197;  #10 
a = 8'd174; b = 8'd198;  #10 
a = 8'd174; b = 8'd199;  #10 
a = 8'd174; b = 8'd200;  #10 
a = 8'd174; b = 8'd201;  #10 
a = 8'd174; b = 8'd202;  #10 
a = 8'd174; b = 8'd203;  #10 
a = 8'd174; b = 8'd204;  #10 
a = 8'd174; b = 8'd205;  #10 
a = 8'd174; b = 8'd206;  #10 
a = 8'd174; b = 8'd207;  #10 
a = 8'd174; b = 8'd208;  #10 
a = 8'd174; b = 8'd209;  #10 
a = 8'd174; b = 8'd210;  #10 
a = 8'd174; b = 8'd211;  #10 
a = 8'd174; b = 8'd212;  #10 
a = 8'd174; b = 8'd213;  #10 
a = 8'd174; b = 8'd214;  #10 
a = 8'd174; b = 8'd215;  #10 
a = 8'd174; b = 8'd216;  #10 
a = 8'd174; b = 8'd217;  #10 
a = 8'd174; b = 8'd218;  #10 
a = 8'd174; b = 8'd219;  #10 
a = 8'd174; b = 8'd220;  #10 
a = 8'd174; b = 8'd221;  #10 
a = 8'd174; b = 8'd222;  #10 
a = 8'd174; b = 8'd223;  #10 
a = 8'd174; b = 8'd224;  #10 
a = 8'd174; b = 8'd225;  #10 
a = 8'd174; b = 8'd226;  #10 
a = 8'd174; b = 8'd227;  #10 
a = 8'd174; b = 8'd228;  #10 
a = 8'd174; b = 8'd229;  #10 
a = 8'd174; b = 8'd230;  #10 
a = 8'd174; b = 8'd231;  #10 
a = 8'd174; b = 8'd232;  #10 
a = 8'd174; b = 8'd233;  #10 
a = 8'd174; b = 8'd234;  #10 
a = 8'd174; b = 8'd235;  #10 
a = 8'd174; b = 8'd236;  #10 
a = 8'd174; b = 8'd237;  #10 
a = 8'd174; b = 8'd238;  #10 
a = 8'd174; b = 8'd239;  #10 
a = 8'd174; b = 8'd240;  #10 
a = 8'd174; b = 8'd241;  #10 
a = 8'd174; b = 8'd242;  #10 
a = 8'd174; b = 8'd243;  #10 
a = 8'd174; b = 8'd244;  #10 
a = 8'd174; b = 8'd245;  #10 
a = 8'd174; b = 8'd246;  #10 
a = 8'd174; b = 8'd247;  #10 
a = 8'd174; b = 8'd248;  #10 
a = 8'd174; b = 8'd249;  #10 
a = 8'd174; b = 8'd250;  #10 
a = 8'd174; b = 8'd251;  #10 
a = 8'd174; b = 8'd252;  #10 
a = 8'd174; b = 8'd253;  #10 
a = 8'd174; b = 8'd254;  #10 
a = 8'd174; b = 8'd255;  #10 
a = 8'd175; b = 8'd0;  #10 
a = 8'd175; b = 8'd1;  #10 
a = 8'd175; b = 8'd2;  #10 
a = 8'd175; b = 8'd3;  #10 
a = 8'd175; b = 8'd4;  #10 
a = 8'd175; b = 8'd5;  #10 
a = 8'd175; b = 8'd6;  #10 
a = 8'd175; b = 8'd7;  #10 
a = 8'd175; b = 8'd8;  #10 
a = 8'd175; b = 8'd9;  #10 
a = 8'd175; b = 8'd10;  #10 
a = 8'd175; b = 8'd11;  #10 
a = 8'd175; b = 8'd12;  #10 
a = 8'd175; b = 8'd13;  #10 
a = 8'd175; b = 8'd14;  #10 
a = 8'd175; b = 8'd15;  #10 
a = 8'd175; b = 8'd16;  #10 
a = 8'd175; b = 8'd17;  #10 
a = 8'd175; b = 8'd18;  #10 
a = 8'd175; b = 8'd19;  #10 
a = 8'd175; b = 8'd20;  #10 
a = 8'd175; b = 8'd21;  #10 
a = 8'd175; b = 8'd22;  #10 
a = 8'd175; b = 8'd23;  #10 
a = 8'd175; b = 8'd24;  #10 
a = 8'd175; b = 8'd25;  #10 
a = 8'd175; b = 8'd26;  #10 
a = 8'd175; b = 8'd27;  #10 
a = 8'd175; b = 8'd28;  #10 
a = 8'd175; b = 8'd29;  #10 
a = 8'd175; b = 8'd30;  #10 
a = 8'd175; b = 8'd31;  #10 
a = 8'd175; b = 8'd32;  #10 
a = 8'd175; b = 8'd33;  #10 
a = 8'd175; b = 8'd34;  #10 
a = 8'd175; b = 8'd35;  #10 
a = 8'd175; b = 8'd36;  #10 
a = 8'd175; b = 8'd37;  #10 
a = 8'd175; b = 8'd38;  #10 
a = 8'd175; b = 8'd39;  #10 
a = 8'd175; b = 8'd40;  #10 
a = 8'd175; b = 8'd41;  #10 
a = 8'd175; b = 8'd42;  #10 
a = 8'd175; b = 8'd43;  #10 
a = 8'd175; b = 8'd44;  #10 
a = 8'd175; b = 8'd45;  #10 
a = 8'd175; b = 8'd46;  #10 
a = 8'd175; b = 8'd47;  #10 
a = 8'd175; b = 8'd48;  #10 
a = 8'd175; b = 8'd49;  #10 
a = 8'd175; b = 8'd50;  #10 
a = 8'd175; b = 8'd51;  #10 
a = 8'd175; b = 8'd52;  #10 
a = 8'd175; b = 8'd53;  #10 
a = 8'd175; b = 8'd54;  #10 
a = 8'd175; b = 8'd55;  #10 
a = 8'd175; b = 8'd56;  #10 
a = 8'd175; b = 8'd57;  #10 
a = 8'd175; b = 8'd58;  #10 
a = 8'd175; b = 8'd59;  #10 
a = 8'd175; b = 8'd60;  #10 
a = 8'd175; b = 8'd61;  #10 
a = 8'd175; b = 8'd62;  #10 
a = 8'd175; b = 8'd63;  #10 
a = 8'd175; b = 8'd64;  #10 
a = 8'd175; b = 8'd65;  #10 
a = 8'd175; b = 8'd66;  #10 
a = 8'd175; b = 8'd67;  #10 
a = 8'd175; b = 8'd68;  #10 
a = 8'd175; b = 8'd69;  #10 
a = 8'd175; b = 8'd70;  #10 
a = 8'd175; b = 8'd71;  #10 
a = 8'd175; b = 8'd72;  #10 
a = 8'd175; b = 8'd73;  #10 
a = 8'd175; b = 8'd74;  #10 
a = 8'd175; b = 8'd75;  #10 
a = 8'd175; b = 8'd76;  #10 
a = 8'd175; b = 8'd77;  #10 
a = 8'd175; b = 8'd78;  #10 
a = 8'd175; b = 8'd79;  #10 
a = 8'd175; b = 8'd80;  #10 
a = 8'd175; b = 8'd81;  #10 
a = 8'd175; b = 8'd82;  #10 
a = 8'd175; b = 8'd83;  #10 
a = 8'd175; b = 8'd84;  #10 
a = 8'd175; b = 8'd85;  #10 
a = 8'd175; b = 8'd86;  #10 
a = 8'd175; b = 8'd87;  #10 
a = 8'd175; b = 8'd88;  #10 
a = 8'd175; b = 8'd89;  #10 
a = 8'd175; b = 8'd90;  #10 
a = 8'd175; b = 8'd91;  #10 
a = 8'd175; b = 8'd92;  #10 
a = 8'd175; b = 8'd93;  #10 
a = 8'd175; b = 8'd94;  #10 
a = 8'd175; b = 8'd95;  #10 
a = 8'd175; b = 8'd96;  #10 
a = 8'd175; b = 8'd97;  #10 
a = 8'd175; b = 8'd98;  #10 
a = 8'd175; b = 8'd99;  #10 
a = 8'd175; b = 8'd100;  #10 
a = 8'd175; b = 8'd101;  #10 
a = 8'd175; b = 8'd102;  #10 
a = 8'd175; b = 8'd103;  #10 
a = 8'd175; b = 8'd104;  #10 
a = 8'd175; b = 8'd105;  #10 
a = 8'd175; b = 8'd106;  #10 
a = 8'd175; b = 8'd107;  #10 
a = 8'd175; b = 8'd108;  #10 
a = 8'd175; b = 8'd109;  #10 
a = 8'd175; b = 8'd110;  #10 
a = 8'd175; b = 8'd111;  #10 
a = 8'd175; b = 8'd112;  #10 
a = 8'd175; b = 8'd113;  #10 
a = 8'd175; b = 8'd114;  #10 
a = 8'd175; b = 8'd115;  #10 
a = 8'd175; b = 8'd116;  #10 
a = 8'd175; b = 8'd117;  #10 
a = 8'd175; b = 8'd118;  #10 
a = 8'd175; b = 8'd119;  #10 
a = 8'd175; b = 8'd120;  #10 
a = 8'd175; b = 8'd121;  #10 
a = 8'd175; b = 8'd122;  #10 
a = 8'd175; b = 8'd123;  #10 
a = 8'd175; b = 8'd124;  #10 
a = 8'd175; b = 8'd125;  #10 
a = 8'd175; b = 8'd126;  #10 
a = 8'd175; b = 8'd127;  #10 
a = 8'd175; b = 8'd128;  #10 
a = 8'd175; b = 8'd129;  #10 
a = 8'd175; b = 8'd130;  #10 
a = 8'd175; b = 8'd131;  #10 
a = 8'd175; b = 8'd132;  #10 
a = 8'd175; b = 8'd133;  #10 
a = 8'd175; b = 8'd134;  #10 
a = 8'd175; b = 8'd135;  #10 
a = 8'd175; b = 8'd136;  #10 
a = 8'd175; b = 8'd137;  #10 
a = 8'd175; b = 8'd138;  #10 
a = 8'd175; b = 8'd139;  #10 
a = 8'd175; b = 8'd140;  #10 
a = 8'd175; b = 8'd141;  #10 
a = 8'd175; b = 8'd142;  #10 
a = 8'd175; b = 8'd143;  #10 
a = 8'd175; b = 8'd144;  #10 
a = 8'd175; b = 8'd145;  #10 
a = 8'd175; b = 8'd146;  #10 
a = 8'd175; b = 8'd147;  #10 
a = 8'd175; b = 8'd148;  #10 
a = 8'd175; b = 8'd149;  #10 
a = 8'd175; b = 8'd150;  #10 
a = 8'd175; b = 8'd151;  #10 
a = 8'd175; b = 8'd152;  #10 
a = 8'd175; b = 8'd153;  #10 
a = 8'd175; b = 8'd154;  #10 
a = 8'd175; b = 8'd155;  #10 
a = 8'd175; b = 8'd156;  #10 
a = 8'd175; b = 8'd157;  #10 
a = 8'd175; b = 8'd158;  #10 
a = 8'd175; b = 8'd159;  #10 
a = 8'd175; b = 8'd160;  #10 
a = 8'd175; b = 8'd161;  #10 
a = 8'd175; b = 8'd162;  #10 
a = 8'd175; b = 8'd163;  #10 
a = 8'd175; b = 8'd164;  #10 
a = 8'd175; b = 8'd165;  #10 
a = 8'd175; b = 8'd166;  #10 
a = 8'd175; b = 8'd167;  #10 
a = 8'd175; b = 8'd168;  #10 
a = 8'd175; b = 8'd169;  #10 
a = 8'd175; b = 8'd170;  #10 
a = 8'd175; b = 8'd171;  #10 
a = 8'd175; b = 8'd172;  #10 
a = 8'd175; b = 8'd173;  #10 
a = 8'd175; b = 8'd174;  #10 
a = 8'd175; b = 8'd175;  #10 
a = 8'd175; b = 8'd176;  #10 
a = 8'd175; b = 8'd177;  #10 
a = 8'd175; b = 8'd178;  #10 
a = 8'd175; b = 8'd179;  #10 
a = 8'd175; b = 8'd180;  #10 
a = 8'd175; b = 8'd181;  #10 
a = 8'd175; b = 8'd182;  #10 
a = 8'd175; b = 8'd183;  #10 
a = 8'd175; b = 8'd184;  #10 
a = 8'd175; b = 8'd185;  #10 
a = 8'd175; b = 8'd186;  #10 
a = 8'd175; b = 8'd187;  #10 
a = 8'd175; b = 8'd188;  #10 
a = 8'd175; b = 8'd189;  #10 
a = 8'd175; b = 8'd190;  #10 
a = 8'd175; b = 8'd191;  #10 
a = 8'd175; b = 8'd192;  #10 
a = 8'd175; b = 8'd193;  #10 
a = 8'd175; b = 8'd194;  #10 
a = 8'd175; b = 8'd195;  #10 
a = 8'd175; b = 8'd196;  #10 
a = 8'd175; b = 8'd197;  #10 
a = 8'd175; b = 8'd198;  #10 
a = 8'd175; b = 8'd199;  #10 
a = 8'd175; b = 8'd200;  #10 
a = 8'd175; b = 8'd201;  #10 
a = 8'd175; b = 8'd202;  #10 
a = 8'd175; b = 8'd203;  #10 
a = 8'd175; b = 8'd204;  #10 
a = 8'd175; b = 8'd205;  #10 
a = 8'd175; b = 8'd206;  #10 
a = 8'd175; b = 8'd207;  #10 
a = 8'd175; b = 8'd208;  #10 
a = 8'd175; b = 8'd209;  #10 
a = 8'd175; b = 8'd210;  #10 
a = 8'd175; b = 8'd211;  #10 
a = 8'd175; b = 8'd212;  #10 
a = 8'd175; b = 8'd213;  #10 
a = 8'd175; b = 8'd214;  #10 
a = 8'd175; b = 8'd215;  #10 
a = 8'd175; b = 8'd216;  #10 
a = 8'd175; b = 8'd217;  #10 
a = 8'd175; b = 8'd218;  #10 
a = 8'd175; b = 8'd219;  #10 
a = 8'd175; b = 8'd220;  #10 
a = 8'd175; b = 8'd221;  #10 
a = 8'd175; b = 8'd222;  #10 
a = 8'd175; b = 8'd223;  #10 
a = 8'd175; b = 8'd224;  #10 
a = 8'd175; b = 8'd225;  #10 
a = 8'd175; b = 8'd226;  #10 
a = 8'd175; b = 8'd227;  #10 
a = 8'd175; b = 8'd228;  #10 
a = 8'd175; b = 8'd229;  #10 
a = 8'd175; b = 8'd230;  #10 
a = 8'd175; b = 8'd231;  #10 
a = 8'd175; b = 8'd232;  #10 
a = 8'd175; b = 8'd233;  #10 
a = 8'd175; b = 8'd234;  #10 
a = 8'd175; b = 8'd235;  #10 
a = 8'd175; b = 8'd236;  #10 
a = 8'd175; b = 8'd237;  #10 
a = 8'd175; b = 8'd238;  #10 
a = 8'd175; b = 8'd239;  #10 
a = 8'd175; b = 8'd240;  #10 
a = 8'd175; b = 8'd241;  #10 
a = 8'd175; b = 8'd242;  #10 
a = 8'd175; b = 8'd243;  #10 
a = 8'd175; b = 8'd244;  #10 
a = 8'd175; b = 8'd245;  #10 
a = 8'd175; b = 8'd246;  #10 
a = 8'd175; b = 8'd247;  #10 
a = 8'd175; b = 8'd248;  #10 
a = 8'd175; b = 8'd249;  #10 
a = 8'd175; b = 8'd250;  #10 
a = 8'd175; b = 8'd251;  #10 
a = 8'd175; b = 8'd252;  #10 
a = 8'd175; b = 8'd253;  #10 
a = 8'd175; b = 8'd254;  #10 
a = 8'd175; b = 8'd255;  #10 
a = 8'd176; b = 8'd0;  #10 
a = 8'd176; b = 8'd1;  #10 
a = 8'd176; b = 8'd2;  #10 
a = 8'd176; b = 8'd3;  #10 
a = 8'd176; b = 8'd4;  #10 
a = 8'd176; b = 8'd5;  #10 
a = 8'd176; b = 8'd6;  #10 
a = 8'd176; b = 8'd7;  #10 
a = 8'd176; b = 8'd8;  #10 
a = 8'd176; b = 8'd9;  #10 
a = 8'd176; b = 8'd10;  #10 
a = 8'd176; b = 8'd11;  #10 
a = 8'd176; b = 8'd12;  #10 
a = 8'd176; b = 8'd13;  #10 
a = 8'd176; b = 8'd14;  #10 
a = 8'd176; b = 8'd15;  #10 
a = 8'd176; b = 8'd16;  #10 
a = 8'd176; b = 8'd17;  #10 
a = 8'd176; b = 8'd18;  #10 
a = 8'd176; b = 8'd19;  #10 
a = 8'd176; b = 8'd20;  #10 
a = 8'd176; b = 8'd21;  #10 
a = 8'd176; b = 8'd22;  #10 
a = 8'd176; b = 8'd23;  #10 
a = 8'd176; b = 8'd24;  #10 
a = 8'd176; b = 8'd25;  #10 
a = 8'd176; b = 8'd26;  #10 
a = 8'd176; b = 8'd27;  #10 
a = 8'd176; b = 8'd28;  #10 
a = 8'd176; b = 8'd29;  #10 
a = 8'd176; b = 8'd30;  #10 
a = 8'd176; b = 8'd31;  #10 
a = 8'd176; b = 8'd32;  #10 
a = 8'd176; b = 8'd33;  #10 
a = 8'd176; b = 8'd34;  #10 
a = 8'd176; b = 8'd35;  #10 
a = 8'd176; b = 8'd36;  #10 
a = 8'd176; b = 8'd37;  #10 
a = 8'd176; b = 8'd38;  #10 
a = 8'd176; b = 8'd39;  #10 
a = 8'd176; b = 8'd40;  #10 
a = 8'd176; b = 8'd41;  #10 
a = 8'd176; b = 8'd42;  #10 
a = 8'd176; b = 8'd43;  #10 
a = 8'd176; b = 8'd44;  #10 
a = 8'd176; b = 8'd45;  #10 
a = 8'd176; b = 8'd46;  #10 
a = 8'd176; b = 8'd47;  #10 
a = 8'd176; b = 8'd48;  #10 
a = 8'd176; b = 8'd49;  #10 
a = 8'd176; b = 8'd50;  #10 
a = 8'd176; b = 8'd51;  #10 
a = 8'd176; b = 8'd52;  #10 
a = 8'd176; b = 8'd53;  #10 
a = 8'd176; b = 8'd54;  #10 
a = 8'd176; b = 8'd55;  #10 
a = 8'd176; b = 8'd56;  #10 
a = 8'd176; b = 8'd57;  #10 
a = 8'd176; b = 8'd58;  #10 
a = 8'd176; b = 8'd59;  #10 
a = 8'd176; b = 8'd60;  #10 
a = 8'd176; b = 8'd61;  #10 
a = 8'd176; b = 8'd62;  #10 
a = 8'd176; b = 8'd63;  #10 
a = 8'd176; b = 8'd64;  #10 
a = 8'd176; b = 8'd65;  #10 
a = 8'd176; b = 8'd66;  #10 
a = 8'd176; b = 8'd67;  #10 
a = 8'd176; b = 8'd68;  #10 
a = 8'd176; b = 8'd69;  #10 
a = 8'd176; b = 8'd70;  #10 
a = 8'd176; b = 8'd71;  #10 
a = 8'd176; b = 8'd72;  #10 
a = 8'd176; b = 8'd73;  #10 
a = 8'd176; b = 8'd74;  #10 
a = 8'd176; b = 8'd75;  #10 
a = 8'd176; b = 8'd76;  #10 
a = 8'd176; b = 8'd77;  #10 
a = 8'd176; b = 8'd78;  #10 
a = 8'd176; b = 8'd79;  #10 
a = 8'd176; b = 8'd80;  #10 
a = 8'd176; b = 8'd81;  #10 
a = 8'd176; b = 8'd82;  #10 
a = 8'd176; b = 8'd83;  #10 
a = 8'd176; b = 8'd84;  #10 
a = 8'd176; b = 8'd85;  #10 
a = 8'd176; b = 8'd86;  #10 
a = 8'd176; b = 8'd87;  #10 
a = 8'd176; b = 8'd88;  #10 
a = 8'd176; b = 8'd89;  #10 
a = 8'd176; b = 8'd90;  #10 
a = 8'd176; b = 8'd91;  #10 
a = 8'd176; b = 8'd92;  #10 
a = 8'd176; b = 8'd93;  #10 
a = 8'd176; b = 8'd94;  #10 
a = 8'd176; b = 8'd95;  #10 
a = 8'd176; b = 8'd96;  #10 
a = 8'd176; b = 8'd97;  #10 
a = 8'd176; b = 8'd98;  #10 
a = 8'd176; b = 8'd99;  #10 
a = 8'd176; b = 8'd100;  #10 
a = 8'd176; b = 8'd101;  #10 
a = 8'd176; b = 8'd102;  #10 
a = 8'd176; b = 8'd103;  #10 
a = 8'd176; b = 8'd104;  #10 
a = 8'd176; b = 8'd105;  #10 
a = 8'd176; b = 8'd106;  #10 
a = 8'd176; b = 8'd107;  #10 
a = 8'd176; b = 8'd108;  #10 
a = 8'd176; b = 8'd109;  #10 
a = 8'd176; b = 8'd110;  #10 
a = 8'd176; b = 8'd111;  #10 
a = 8'd176; b = 8'd112;  #10 
a = 8'd176; b = 8'd113;  #10 
a = 8'd176; b = 8'd114;  #10 
a = 8'd176; b = 8'd115;  #10 
a = 8'd176; b = 8'd116;  #10 
a = 8'd176; b = 8'd117;  #10 
a = 8'd176; b = 8'd118;  #10 
a = 8'd176; b = 8'd119;  #10 
a = 8'd176; b = 8'd120;  #10 
a = 8'd176; b = 8'd121;  #10 
a = 8'd176; b = 8'd122;  #10 
a = 8'd176; b = 8'd123;  #10 
a = 8'd176; b = 8'd124;  #10 
a = 8'd176; b = 8'd125;  #10 
a = 8'd176; b = 8'd126;  #10 
a = 8'd176; b = 8'd127;  #10 
a = 8'd176; b = 8'd128;  #10 
a = 8'd176; b = 8'd129;  #10 
a = 8'd176; b = 8'd130;  #10 
a = 8'd176; b = 8'd131;  #10 
a = 8'd176; b = 8'd132;  #10 
a = 8'd176; b = 8'd133;  #10 
a = 8'd176; b = 8'd134;  #10 
a = 8'd176; b = 8'd135;  #10 
a = 8'd176; b = 8'd136;  #10 
a = 8'd176; b = 8'd137;  #10 
a = 8'd176; b = 8'd138;  #10 
a = 8'd176; b = 8'd139;  #10 
a = 8'd176; b = 8'd140;  #10 
a = 8'd176; b = 8'd141;  #10 
a = 8'd176; b = 8'd142;  #10 
a = 8'd176; b = 8'd143;  #10 
a = 8'd176; b = 8'd144;  #10 
a = 8'd176; b = 8'd145;  #10 
a = 8'd176; b = 8'd146;  #10 
a = 8'd176; b = 8'd147;  #10 
a = 8'd176; b = 8'd148;  #10 
a = 8'd176; b = 8'd149;  #10 
a = 8'd176; b = 8'd150;  #10 
a = 8'd176; b = 8'd151;  #10 
a = 8'd176; b = 8'd152;  #10 
a = 8'd176; b = 8'd153;  #10 
a = 8'd176; b = 8'd154;  #10 
a = 8'd176; b = 8'd155;  #10 
a = 8'd176; b = 8'd156;  #10 
a = 8'd176; b = 8'd157;  #10 
a = 8'd176; b = 8'd158;  #10 
a = 8'd176; b = 8'd159;  #10 
a = 8'd176; b = 8'd160;  #10 
a = 8'd176; b = 8'd161;  #10 
a = 8'd176; b = 8'd162;  #10 
a = 8'd176; b = 8'd163;  #10 
a = 8'd176; b = 8'd164;  #10 
a = 8'd176; b = 8'd165;  #10 
a = 8'd176; b = 8'd166;  #10 
a = 8'd176; b = 8'd167;  #10 
a = 8'd176; b = 8'd168;  #10 
a = 8'd176; b = 8'd169;  #10 
a = 8'd176; b = 8'd170;  #10 
a = 8'd176; b = 8'd171;  #10 
a = 8'd176; b = 8'd172;  #10 
a = 8'd176; b = 8'd173;  #10 
a = 8'd176; b = 8'd174;  #10 
a = 8'd176; b = 8'd175;  #10 
a = 8'd176; b = 8'd176;  #10 
a = 8'd176; b = 8'd177;  #10 
a = 8'd176; b = 8'd178;  #10 
a = 8'd176; b = 8'd179;  #10 
a = 8'd176; b = 8'd180;  #10 
a = 8'd176; b = 8'd181;  #10 
a = 8'd176; b = 8'd182;  #10 
a = 8'd176; b = 8'd183;  #10 
a = 8'd176; b = 8'd184;  #10 
a = 8'd176; b = 8'd185;  #10 
a = 8'd176; b = 8'd186;  #10 
a = 8'd176; b = 8'd187;  #10 
a = 8'd176; b = 8'd188;  #10 
a = 8'd176; b = 8'd189;  #10 
a = 8'd176; b = 8'd190;  #10 
a = 8'd176; b = 8'd191;  #10 
a = 8'd176; b = 8'd192;  #10 
a = 8'd176; b = 8'd193;  #10 
a = 8'd176; b = 8'd194;  #10 
a = 8'd176; b = 8'd195;  #10 
a = 8'd176; b = 8'd196;  #10 
a = 8'd176; b = 8'd197;  #10 
a = 8'd176; b = 8'd198;  #10 
a = 8'd176; b = 8'd199;  #10 
a = 8'd176; b = 8'd200;  #10 
a = 8'd176; b = 8'd201;  #10 
a = 8'd176; b = 8'd202;  #10 
a = 8'd176; b = 8'd203;  #10 
a = 8'd176; b = 8'd204;  #10 
a = 8'd176; b = 8'd205;  #10 
a = 8'd176; b = 8'd206;  #10 
a = 8'd176; b = 8'd207;  #10 
a = 8'd176; b = 8'd208;  #10 
a = 8'd176; b = 8'd209;  #10 
a = 8'd176; b = 8'd210;  #10 
a = 8'd176; b = 8'd211;  #10 
a = 8'd176; b = 8'd212;  #10 
a = 8'd176; b = 8'd213;  #10 
a = 8'd176; b = 8'd214;  #10 
a = 8'd176; b = 8'd215;  #10 
a = 8'd176; b = 8'd216;  #10 
a = 8'd176; b = 8'd217;  #10 
a = 8'd176; b = 8'd218;  #10 
a = 8'd176; b = 8'd219;  #10 
a = 8'd176; b = 8'd220;  #10 
a = 8'd176; b = 8'd221;  #10 
a = 8'd176; b = 8'd222;  #10 
a = 8'd176; b = 8'd223;  #10 
a = 8'd176; b = 8'd224;  #10 
a = 8'd176; b = 8'd225;  #10 
a = 8'd176; b = 8'd226;  #10 
a = 8'd176; b = 8'd227;  #10 
a = 8'd176; b = 8'd228;  #10 
a = 8'd176; b = 8'd229;  #10 
a = 8'd176; b = 8'd230;  #10 
a = 8'd176; b = 8'd231;  #10 
a = 8'd176; b = 8'd232;  #10 
a = 8'd176; b = 8'd233;  #10 
a = 8'd176; b = 8'd234;  #10 
a = 8'd176; b = 8'd235;  #10 
a = 8'd176; b = 8'd236;  #10 
a = 8'd176; b = 8'd237;  #10 
a = 8'd176; b = 8'd238;  #10 
a = 8'd176; b = 8'd239;  #10 
a = 8'd176; b = 8'd240;  #10 
a = 8'd176; b = 8'd241;  #10 
a = 8'd176; b = 8'd242;  #10 
a = 8'd176; b = 8'd243;  #10 
a = 8'd176; b = 8'd244;  #10 
a = 8'd176; b = 8'd245;  #10 
a = 8'd176; b = 8'd246;  #10 
a = 8'd176; b = 8'd247;  #10 
a = 8'd176; b = 8'd248;  #10 
a = 8'd176; b = 8'd249;  #10 
a = 8'd176; b = 8'd250;  #10 
a = 8'd176; b = 8'd251;  #10 
a = 8'd176; b = 8'd252;  #10 
a = 8'd176; b = 8'd253;  #10 
a = 8'd176; b = 8'd254;  #10 
a = 8'd176; b = 8'd255;  #10 
a = 8'd177; b = 8'd0;  #10 
a = 8'd177; b = 8'd1;  #10 
a = 8'd177; b = 8'd2;  #10 
a = 8'd177; b = 8'd3;  #10 
a = 8'd177; b = 8'd4;  #10 
a = 8'd177; b = 8'd5;  #10 
a = 8'd177; b = 8'd6;  #10 
a = 8'd177; b = 8'd7;  #10 
a = 8'd177; b = 8'd8;  #10 
a = 8'd177; b = 8'd9;  #10 
a = 8'd177; b = 8'd10;  #10 
a = 8'd177; b = 8'd11;  #10 
a = 8'd177; b = 8'd12;  #10 
a = 8'd177; b = 8'd13;  #10 
a = 8'd177; b = 8'd14;  #10 
a = 8'd177; b = 8'd15;  #10 
a = 8'd177; b = 8'd16;  #10 
a = 8'd177; b = 8'd17;  #10 
a = 8'd177; b = 8'd18;  #10 
a = 8'd177; b = 8'd19;  #10 
a = 8'd177; b = 8'd20;  #10 
a = 8'd177; b = 8'd21;  #10 
a = 8'd177; b = 8'd22;  #10 
a = 8'd177; b = 8'd23;  #10 
a = 8'd177; b = 8'd24;  #10 
a = 8'd177; b = 8'd25;  #10 
a = 8'd177; b = 8'd26;  #10 
a = 8'd177; b = 8'd27;  #10 
a = 8'd177; b = 8'd28;  #10 
a = 8'd177; b = 8'd29;  #10 
a = 8'd177; b = 8'd30;  #10 
a = 8'd177; b = 8'd31;  #10 
a = 8'd177; b = 8'd32;  #10 
a = 8'd177; b = 8'd33;  #10 
a = 8'd177; b = 8'd34;  #10 
a = 8'd177; b = 8'd35;  #10 
a = 8'd177; b = 8'd36;  #10 
a = 8'd177; b = 8'd37;  #10 
a = 8'd177; b = 8'd38;  #10 
a = 8'd177; b = 8'd39;  #10 
a = 8'd177; b = 8'd40;  #10 
a = 8'd177; b = 8'd41;  #10 
a = 8'd177; b = 8'd42;  #10 
a = 8'd177; b = 8'd43;  #10 
a = 8'd177; b = 8'd44;  #10 
a = 8'd177; b = 8'd45;  #10 
a = 8'd177; b = 8'd46;  #10 
a = 8'd177; b = 8'd47;  #10 
a = 8'd177; b = 8'd48;  #10 
a = 8'd177; b = 8'd49;  #10 
a = 8'd177; b = 8'd50;  #10 
a = 8'd177; b = 8'd51;  #10 
a = 8'd177; b = 8'd52;  #10 
a = 8'd177; b = 8'd53;  #10 
a = 8'd177; b = 8'd54;  #10 
a = 8'd177; b = 8'd55;  #10 
a = 8'd177; b = 8'd56;  #10 
a = 8'd177; b = 8'd57;  #10 
a = 8'd177; b = 8'd58;  #10 
a = 8'd177; b = 8'd59;  #10 
a = 8'd177; b = 8'd60;  #10 
a = 8'd177; b = 8'd61;  #10 
a = 8'd177; b = 8'd62;  #10 
a = 8'd177; b = 8'd63;  #10 
a = 8'd177; b = 8'd64;  #10 
a = 8'd177; b = 8'd65;  #10 
a = 8'd177; b = 8'd66;  #10 
a = 8'd177; b = 8'd67;  #10 
a = 8'd177; b = 8'd68;  #10 
a = 8'd177; b = 8'd69;  #10 
a = 8'd177; b = 8'd70;  #10 
a = 8'd177; b = 8'd71;  #10 
a = 8'd177; b = 8'd72;  #10 
a = 8'd177; b = 8'd73;  #10 
a = 8'd177; b = 8'd74;  #10 
a = 8'd177; b = 8'd75;  #10 
a = 8'd177; b = 8'd76;  #10 
a = 8'd177; b = 8'd77;  #10 
a = 8'd177; b = 8'd78;  #10 
a = 8'd177; b = 8'd79;  #10 
a = 8'd177; b = 8'd80;  #10 
a = 8'd177; b = 8'd81;  #10 
a = 8'd177; b = 8'd82;  #10 
a = 8'd177; b = 8'd83;  #10 
a = 8'd177; b = 8'd84;  #10 
a = 8'd177; b = 8'd85;  #10 
a = 8'd177; b = 8'd86;  #10 
a = 8'd177; b = 8'd87;  #10 
a = 8'd177; b = 8'd88;  #10 
a = 8'd177; b = 8'd89;  #10 
a = 8'd177; b = 8'd90;  #10 
a = 8'd177; b = 8'd91;  #10 
a = 8'd177; b = 8'd92;  #10 
a = 8'd177; b = 8'd93;  #10 
a = 8'd177; b = 8'd94;  #10 
a = 8'd177; b = 8'd95;  #10 
a = 8'd177; b = 8'd96;  #10 
a = 8'd177; b = 8'd97;  #10 
a = 8'd177; b = 8'd98;  #10 
a = 8'd177; b = 8'd99;  #10 
a = 8'd177; b = 8'd100;  #10 
a = 8'd177; b = 8'd101;  #10 
a = 8'd177; b = 8'd102;  #10 
a = 8'd177; b = 8'd103;  #10 
a = 8'd177; b = 8'd104;  #10 
a = 8'd177; b = 8'd105;  #10 
a = 8'd177; b = 8'd106;  #10 
a = 8'd177; b = 8'd107;  #10 
a = 8'd177; b = 8'd108;  #10 
a = 8'd177; b = 8'd109;  #10 
a = 8'd177; b = 8'd110;  #10 
a = 8'd177; b = 8'd111;  #10 
a = 8'd177; b = 8'd112;  #10 
a = 8'd177; b = 8'd113;  #10 
a = 8'd177; b = 8'd114;  #10 
a = 8'd177; b = 8'd115;  #10 
a = 8'd177; b = 8'd116;  #10 
a = 8'd177; b = 8'd117;  #10 
a = 8'd177; b = 8'd118;  #10 
a = 8'd177; b = 8'd119;  #10 
a = 8'd177; b = 8'd120;  #10 
a = 8'd177; b = 8'd121;  #10 
a = 8'd177; b = 8'd122;  #10 
a = 8'd177; b = 8'd123;  #10 
a = 8'd177; b = 8'd124;  #10 
a = 8'd177; b = 8'd125;  #10 
a = 8'd177; b = 8'd126;  #10 
a = 8'd177; b = 8'd127;  #10 
a = 8'd177; b = 8'd128;  #10 
a = 8'd177; b = 8'd129;  #10 
a = 8'd177; b = 8'd130;  #10 
a = 8'd177; b = 8'd131;  #10 
a = 8'd177; b = 8'd132;  #10 
a = 8'd177; b = 8'd133;  #10 
a = 8'd177; b = 8'd134;  #10 
a = 8'd177; b = 8'd135;  #10 
a = 8'd177; b = 8'd136;  #10 
a = 8'd177; b = 8'd137;  #10 
a = 8'd177; b = 8'd138;  #10 
a = 8'd177; b = 8'd139;  #10 
a = 8'd177; b = 8'd140;  #10 
a = 8'd177; b = 8'd141;  #10 
a = 8'd177; b = 8'd142;  #10 
a = 8'd177; b = 8'd143;  #10 
a = 8'd177; b = 8'd144;  #10 
a = 8'd177; b = 8'd145;  #10 
a = 8'd177; b = 8'd146;  #10 
a = 8'd177; b = 8'd147;  #10 
a = 8'd177; b = 8'd148;  #10 
a = 8'd177; b = 8'd149;  #10 
a = 8'd177; b = 8'd150;  #10 
a = 8'd177; b = 8'd151;  #10 
a = 8'd177; b = 8'd152;  #10 
a = 8'd177; b = 8'd153;  #10 
a = 8'd177; b = 8'd154;  #10 
a = 8'd177; b = 8'd155;  #10 
a = 8'd177; b = 8'd156;  #10 
a = 8'd177; b = 8'd157;  #10 
a = 8'd177; b = 8'd158;  #10 
a = 8'd177; b = 8'd159;  #10 
a = 8'd177; b = 8'd160;  #10 
a = 8'd177; b = 8'd161;  #10 
a = 8'd177; b = 8'd162;  #10 
a = 8'd177; b = 8'd163;  #10 
a = 8'd177; b = 8'd164;  #10 
a = 8'd177; b = 8'd165;  #10 
a = 8'd177; b = 8'd166;  #10 
a = 8'd177; b = 8'd167;  #10 
a = 8'd177; b = 8'd168;  #10 
a = 8'd177; b = 8'd169;  #10 
a = 8'd177; b = 8'd170;  #10 
a = 8'd177; b = 8'd171;  #10 
a = 8'd177; b = 8'd172;  #10 
a = 8'd177; b = 8'd173;  #10 
a = 8'd177; b = 8'd174;  #10 
a = 8'd177; b = 8'd175;  #10 
a = 8'd177; b = 8'd176;  #10 
a = 8'd177; b = 8'd177;  #10 
a = 8'd177; b = 8'd178;  #10 
a = 8'd177; b = 8'd179;  #10 
a = 8'd177; b = 8'd180;  #10 
a = 8'd177; b = 8'd181;  #10 
a = 8'd177; b = 8'd182;  #10 
a = 8'd177; b = 8'd183;  #10 
a = 8'd177; b = 8'd184;  #10 
a = 8'd177; b = 8'd185;  #10 
a = 8'd177; b = 8'd186;  #10 
a = 8'd177; b = 8'd187;  #10 
a = 8'd177; b = 8'd188;  #10 
a = 8'd177; b = 8'd189;  #10 
a = 8'd177; b = 8'd190;  #10 
a = 8'd177; b = 8'd191;  #10 
a = 8'd177; b = 8'd192;  #10 
a = 8'd177; b = 8'd193;  #10 
a = 8'd177; b = 8'd194;  #10 
a = 8'd177; b = 8'd195;  #10 
a = 8'd177; b = 8'd196;  #10 
a = 8'd177; b = 8'd197;  #10 
a = 8'd177; b = 8'd198;  #10 
a = 8'd177; b = 8'd199;  #10 
a = 8'd177; b = 8'd200;  #10 
a = 8'd177; b = 8'd201;  #10 
a = 8'd177; b = 8'd202;  #10 
a = 8'd177; b = 8'd203;  #10 
a = 8'd177; b = 8'd204;  #10 
a = 8'd177; b = 8'd205;  #10 
a = 8'd177; b = 8'd206;  #10 
a = 8'd177; b = 8'd207;  #10 
a = 8'd177; b = 8'd208;  #10 
a = 8'd177; b = 8'd209;  #10 
a = 8'd177; b = 8'd210;  #10 
a = 8'd177; b = 8'd211;  #10 
a = 8'd177; b = 8'd212;  #10 
a = 8'd177; b = 8'd213;  #10 
a = 8'd177; b = 8'd214;  #10 
a = 8'd177; b = 8'd215;  #10 
a = 8'd177; b = 8'd216;  #10 
a = 8'd177; b = 8'd217;  #10 
a = 8'd177; b = 8'd218;  #10 
a = 8'd177; b = 8'd219;  #10 
a = 8'd177; b = 8'd220;  #10 
a = 8'd177; b = 8'd221;  #10 
a = 8'd177; b = 8'd222;  #10 
a = 8'd177; b = 8'd223;  #10 
a = 8'd177; b = 8'd224;  #10 
a = 8'd177; b = 8'd225;  #10 
a = 8'd177; b = 8'd226;  #10 
a = 8'd177; b = 8'd227;  #10 
a = 8'd177; b = 8'd228;  #10 
a = 8'd177; b = 8'd229;  #10 
a = 8'd177; b = 8'd230;  #10 
a = 8'd177; b = 8'd231;  #10 
a = 8'd177; b = 8'd232;  #10 
a = 8'd177; b = 8'd233;  #10 
a = 8'd177; b = 8'd234;  #10 
a = 8'd177; b = 8'd235;  #10 
a = 8'd177; b = 8'd236;  #10 
a = 8'd177; b = 8'd237;  #10 
a = 8'd177; b = 8'd238;  #10 
a = 8'd177; b = 8'd239;  #10 
a = 8'd177; b = 8'd240;  #10 
a = 8'd177; b = 8'd241;  #10 
a = 8'd177; b = 8'd242;  #10 
a = 8'd177; b = 8'd243;  #10 
a = 8'd177; b = 8'd244;  #10 
a = 8'd177; b = 8'd245;  #10 
a = 8'd177; b = 8'd246;  #10 
a = 8'd177; b = 8'd247;  #10 
a = 8'd177; b = 8'd248;  #10 
a = 8'd177; b = 8'd249;  #10 
a = 8'd177; b = 8'd250;  #10 
a = 8'd177; b = 8'd251;  #10 
a = 8'd177; b = 8'd252;  #10 
a = 8'd177; b = 8'd253;  #10 
a = 8'd177; b = 8'd254;  #10 
a = 8'd177; b = 8'd255;  #10 
a = 8'd178; b = 8'd0;  #10 
a = 8'd178; b = 8'd1;  #10 
a = 8'd178; b = 8'd2;  #10 
a = 8'd178; b = 8'd3;  #10 
a = 8'd178; b = 8'd4;  #10 
a = 8'd178; b = 8'd5;  #10 
a = 8'd178; b = 8'd6;  #10 
a = 8'd178; b = 8'd7;  #10 
a = 8'd178; b = 8'd8;  #10 
a = 8'd178; b = 8'd9;  #10 
a = 8'd178; b = 8'd10;  #10 
a = 8'd178; b = 8'd11;  #10 
a = 8'd178; b = 8'd12;  #10 
a = 8'd178; b = 8'd13;  #10 
a = 8'd178; b = 8'd14;  #10 
a = 8'd178; b = 8'd15;  #10 
a = 8'd178; b = 8'd16;  #10 
a = 8'd178; b = 8'd17;  #10 
a = 8'd178; b = 8'd18;  #10 
a = 8'd178; b = 8'd19;  #10 
a = 8'd178; b = 8'd20;  #10 
a = 8'd178; b = 8'd21;  #10 
a = 8'd178; b = 8'd22;  #10 
a = 8'd178; b = 8'd23;  #10 
a = 8'd178; b = 8'd24;  #10 
a = 8'd178; b = 8'd25;  #10 
a = 8'd178; b = 8'd26;  #10 
a = 8'd178; b = 8'd27;  #10 
a = 8'd178; b = 8'd28;  #10 
a = 8'd178; b = 8'd29;  #10 
a = 8'd178; b = 8'd30;  #10 
a = 8'd178; b = 8'd31;  #10 
a = 8'd178; b = 8'd32;  #10 
a = 8'd178; b = 8'd33;  #10 
a = 8'd178; b = 8'd34;  #10 
a = 8'd178; b = 8'd35;  #10 
a = 8'd178; b = 8'd36;  #10 
a = 8'd178; b = 8'd37;  #10 
a = 8'd178; b = 8'd38;  #10 
a = 8'd178; b = 8'd39;  #10 
a = 8'd178; b = 8'd40;  #10 
a = 8'd178; b = 8'd41;  #10 
a = 8'd178; b = 8'd42;  #10 
a = 8'd178; b = 8'd43;  #10 
a = 8'd178; b = 8'd44;  #10 
a = 8'd178; b = 8'd45;  #10 
a = 8'd178; b = 8'd46;  #10 
a = 8'd178; b = 8'd47;  #10 
a = 8'd178; b = 8'd48;  #10 
a = 8'd178; b = 8'd49;  #10 
a = 8'd178; b = 8'd50;  #10 
a = 8'd178; b = 8'd51;  #10 
a = 8'd178; b = 8'd52;  #10 
a = 8'd178; b = 8'd53;  #10 
a = 8'd178; b = 8'd54;  #10 
a = 8'd178; b = 8'd55;  #10 
a = 8'd178; b = 8'd56;  #10 
a = 8'd178; b = 8'd57;  #10 
a = 8'd178; b = 8'd58;  #10 
a = 8'd178; b = 8'd59;  #10 
a = 8'd178; b = 8'd60;  #10 
a = 8'd178; b = 8'd61;  #10 
a = 8'd178; b = 8'd62;  #10 
a = 8'd178; b = 8'd63;  #10 
a = 8'd178; b = 8'd64;  #10 
a = 8'd178; b = 8'd65;  #10 
a = 8'd178; b = 8'd66;  #10 
a = 8'd178; b = 8'd67;  #10 
a = 8'd178; b = 8'd68;  #10 
a = 8'd178; b = 8'd69;  #10 
a = 8'd178; b = 8'd70;  #10 
a = 8'd178; b = 8'd71;  #10 
a = 8'd178; b = 8'd72;  #10 
a = 8'd178; b = 8'd73;  #10 
a = 8'd178; b = 8'd74;  #10 
a = 8'd178; b = 8'd75;  #10 
a = 8'd178; b = 8'd76;  #10 
a = 8'd178; b = 8'd77;  #10 
a = 8'd178; b = 8'd78;  #10 
a = 8'd178; b = 8'd79;  #10 
a = 8'd178; b = 8'd80;  #10 
a = 8'd178; b = 8'd81;  #10 
a = 8'd178; b = 8'd82;  #10 
a = 8'd178; b = 8'd83;  #10 
a = 8'd178; b = 8'd84;  #10 
a = 8'd178; b = 8'd85;  #10 
a = 8'd178; b = 8'd86;  #10 
a = 8'd178; b = 8'd87;  #10 
a = 8'd178; b = 8'd88;  #10 
a = 8'd178; b = 8'd89;  #10 
a = 8'd178; b = 8'd90;  #10 
a = 8'd178; b = 8'd91;  #10 
a = 8'd178; b = 8'd92;  #10 
a = 8'd178; b = 8'd93;  #10 
a = 8'd178; b = 8'd94;  #10 
a = 8'd178; b = 8'd95;  #10 
a = 8'd178; b = 8'd96;  #10 
a = 8'd178; b = 8'd97;  #10 
a = 8'd178; b = 8'd98;  #10 
a = 8'd178; b = 8'd99;  #10 
a = 8'd178; b = 8'd100;  #10 
a = 8'd178; b = 8'd101;  #10 
a = 8'd178; b = 8'd102;  #10 
a = 8'd178; b = 8'd103;  #10 
a = 8'd178; b = 8'd104;  #10 
a = 8'd178; b = 8'd105;  #10 
a = 8'd178; b = 8'd106;  #10 
a = 8'd178; b = 8'd107;  #10 
a = 8'd178; b = 8'd108;  #10 
a = 8'd178; b = 8'd109;  #10 
a = 8'd178; b = 8'd110;  #10 
a = 8'd178; b = 8'd111;  #10 
a = 8'd178; b = 8'd112;  #10 
a = 8'd178; b = 8'd113;  #10 
a = 8'd178; b = 8'd114;  #10 
a = 8'd178; b = 8'd115;  #10 
a = 8'd178; b = 8'd116;  #10 
a = 8'd178; b = 8'd117;  #10 
a = 8'd178; b = 8'd118;  #10 
a = 8'd178; b = 8'd119;  #10 
a = 8'd178; b = 8'd120;  #10 
a = 8'd178; b = 8'd121;  #10 
a = 8'd178; b = 8'd122;  #10 
a = 8'd178; b = 8'd123;  #10 
a = 8'd178; b = 8'd124;  #10 
a = 8'd178; b = 8'd125;  #10 
a = 8'd178; b = 8'd126;  #10 
a = 8'd178; b = 8'd127;  #10 
a = 8'd178; b = 8'd128;  #10 
a = 8'd178; b = 8'd129;  #10 
a = 8'd178; b = 8'd130;  #10 
a = 8'd178; b = 8'd131;  #10 
a = 8'd178; b = 8'd132;  #10 
a = 8'd178; b = 8'd133;  #10 
a = 8'd178; b = 8'd134;  #10 
a = 8'd178; b = 8'd135;  #10 
a = 8'd178; b = 8'd136;  #10 
a = 8'd178; b = 8'd137;  #10 
a = 8'd178; b = 8'd138;  #10 
a = 8'd178; b = 8'd139;  #10 
a = 8'd178; b = 8'd140;  #10 
a = 8'd178; b = 8'd141;  #10 
a = 8'd178; b = 8'd142;  #10 
a = 8'd178; b = 8'd143;  #10 
a = 8'd178; b = 8'd144;  #10 
a = 8'd178; b = 8'd145;  #10 
a = 8'd178; b = 8'd146;  #10 
a = 8'd178; b = 8'd147;  #10 
a = 8'd178; b = 8'd148;  #10 
a = 8'd178; b = 8'd149;  #10 
a = 8'd178; b = 8'd150;  #10 
a = 8'd178; b = 8'd151;  #10 
a = 8'd178; b = 8'd152;  #10 
a = 8'd178; b = 8'd153;  #10 
a = 8'd178; b = 8'd154;  #10 
a = 8'd178; b = 8'd155;  #10 
a = 8'd178; b = 8'd156;  #10 
a = 8'd178; b = 8'd157;  #10 
a = 8'd178; b = 8'd158;  #10 
a = 8'd178; b = 8'd159;  #10 
a = 8'd178; b = 8'd160;  #10 
a = 8'd178; b = 8'd161;  #10 
a = 8'd178; b = 8'd162;  #10 
a = 8'd178; b = 8'd163;  #10 
a = 8'd178; b = 8'd164;  #10 
a = 8'd178; b = 8'd165;  #10 
a = 8'd178; b = 8'd166;  #10 
a = 8'd178; b = 8'd167;  #10 
a = 8'd178; b = 8'd168;  #10 
a = 8'd178; b = 8'd169;  #10 
a = 8'd178; b = 8'd170;  #10 
a = 8'd178; b = 8'd171;  #10 
a = 8'd178; b = 8'd172;  #10 
a = 8'd178; b = 8'd173;  #10 
a = 8'd178; b = 8'd174;  #10 
a = 8'd178; b = 8'd175;  #10 
a = 8'd178; b = 8'd176;  #10 
a = 8'd178; b = 8'd177;  #10 
a = 8'd178; b = 8'd178;  #10 
a = 8'd178; b = 8'd179;  #10 
a = 8'd178; b = 8'd180;  #10 
a = 8'd178; b = 8'd181;  #10 
a = 8'd178; b = 8'd182;  #10 
a = 8'd178; b = 8'd183;  #10 
a = 8'd178; b = 8'd184;  #10 
a = 8'd178; b = 8'd185;  #10 
a = 8'd178; b = 8'd186;  #10 
a = 8'd178; b = 8'd187;  #10 
a = 8'd178; b = 8'd188;  #10 
a = 8'd178; b = 8'd189;  #10 
a = 8'd178; b = 8'd190;  #10 
a = 8'd178; b = 8'd191;  #10 
a = 8'd178; b = 8'd192;  #10 
a = 8'd178; b = 8'd193;  #10 
a = 8'd178; b = 8'd194;  #10 
a = 8'd178; b = 8'd195;  #10 
a = 8'd178; b = 8'd196;  #10 
a = 8'd178; b = 8'd197;  #10 
a = 8'd178; b = 8'd198;  #10 
a = 8'd178; b = 8'd199;  #10 
a = 8'd178; b = 8'd200;  #10 
a = 8'd178; b = 8'd201;  #10 
a = 8'd178; b = 8'd202;  #10 
a = 8'd178; b = 8'd203;  #10 
a = 8'd178; b = 8'd204;  #10 
a = 8'd178; b = 8'd205;  #10 
a = 8'd178; b = 8'd206;  #10 
a = 8'd178; b = 8'd207;  #10 
a = 8'd178; b = 8'd208;  #10 
a = 8'd178; b = 8'd209;  #10 
a = 8'd178; b = 8'd210;  #10 
a = 8'd178; b = 8'd211;  #10 
a = 8'd178; b = 8'd212;  #10 
a = 8'd178; b = 8'd213;  #10 
a = 8'd178; b = 8'd214;  #10 
a = 8'd178; b = 8'd215;  #10 
a = 8'd178; b = 8'd216;  #10 
a = 8'd178; b = 8'd217;  #10 
a = 8'd178; b = 8'd218;  #10 
a = 8'd178; b = 8'd219;  #10 
a = 8'd178; b = 8'd220;  #10 
a = 8'd178; b = 8'd221;  #10 
a = 8'd178; b = 8'd222;  #10 
a = 8'd178; b = 8'd223;  #10 
a = 8'd178; b = 8'd224;  #10 
a = 8'd178; b = 8'd225;  #10 
a = 8'd178; b = 8'd226;  #10 
a = 8'd178; b = 8'd227;  #10 
a = 8'd178; b = 8'd228;  #10 
a = 8'd178; b = 8'd229;  #10 
a = 8'd178; b = 8'd230;  #10 
a = 8'd178; b = 8'd231;  #10 
a = 8'd178; b = 8'd232;  #10 
a = 8'd178; b = 8'd233;  #10 
a = 8'd178; b = 8'd234;  #10 
a = 8'd178; b = 8'd235;  #10 
a = 8'd178; b = 8'd236;  #10 
a = 8'd178; b = 8'd237;  #10 
a = 8'd178; b = 8'd238;  #10 
a = 8'd178; b = 8'd239;  #10 
a = 8'd178; b = 8'd240;  #10 
a = 8'd178; b = 8'd241;  #10 
a = 8'd178; b = 8'd242;  #10 
a = 8'd178; b = 8'd243;  #10 
a = 8'd178; b = 8'd244;  #10 
a = 8'd178; b = 8'd245;  #10 
a = 8'd178; b = 8'd246;  #10 
a = 8'd178; b = 8'd247;  #10 
a = 8'd178; b = 8'd248;  #10 
a = 8'd178; b = 8'd249;  #10 
a = 8'd178; b = 8'd250;  #10 
a = 8'd178; b = 8'd251;  #10 
a = 8'd178; b = 8'd252;  #10 
a = 8'd178; b = 8'd253;  #10 
a = 8'd178; b = 8'd254;  #10 
a = 8'd178; b = 8'd255;  #10 
a = 8'd179; b = 8'd0;  #10 
a = 8'd179; b = 8'd1;  #10 
a = 8'd179; b = 8'd2;  #10 
a = 8'd179; b = 8'd3;  #10 
a = 8'd179; b = 8'd4;  #10 
a = 8'd179; b = 8'd5;  #10 
a = 8'd179; b = 8'd6;  #10 
a = 8'd179; b = 8'd7;  #10 
a = 8'd179; b = 8'd8;  #10 
a = 8'd179; b = 8'd9;  #10 
a = 8'd179; b = 8'd10;  #10 
a = 8'd179; b = 8'd11;  #10 
a = 8'd179; b = 8'd12;  #10 
a = 8'd179; b = 8'd13;  #10 
a = 8'd179; b = 8'd14;  #10 
a = 8'd179; b = 8'd15;  #10 
a = 8'd179; b = 8'd16;  #10 
a = 8'd179; b = 8'd17;  #10 
a = 8'd179; b = 8'd18;  #10 
a = 8'd179; b = 8'd19;  #10 
a = 8'd179; b = 8'd20;  #10 
a = 8'd179; b = 8'd21;  #10 
a = 8'd179; b = 8'd22;  #10 
a = 8'd179; b = 8'd23;  #10 
a = 8'd179; b = 8'd24;  #10 
a = 8'd179; b = 8'd25;  #10 
a = 8'd179; b = 8'd26;  #10 
a = 8'd179; b = 8'd27;  #10 
a = 8'd179; b = 8'd28;  #10 
a = 8'd179; b = 8'd29;  #10 
a = 8'd179; b = 8'd30;  #10 
a = 8'd179; b = 8'd31;  #10 
a = 8'd179; b = 8'd32;  #10 
a = 8'd179; b = 8'd33;  #10 
a = 8'd179; b = 8'd34;  #10 
a = 8'd179; b = 8'd35;  #10 
a = 8'd179; b = 8'd36;  #10 
a = 8'd179; b = 8'd37;  #10 
a = 8'd179; b = 8'd38;  #10 
a = 8'd179; b = 8'd39;  #10 
a = 8'd179; b = 8'd40;  #10 
a = 8'd179; b = 8'd41;  #10 
a = 8'd179; b = 8'd42;  #10 
a = 8'd179; b = 8'd43;  #10 
a = 8'd179; b = 8'd44;  #10 
a = 8'd179; b = 8'd45;  #10 
a = 8'd179; b = 8'd46;  #10 
a = 8'd179; b = 8'd47;  #10 
a = 8'd179; b = 8'd48;  #10 
a = 8'd179; b = 8'd49;  #10 
a = 8'd179; b = 8'd50;  #10 
a = 8'd179; b = 8'd51;  #10 
a = 8'd179; b = 8'd52;  #10 
a = 8'd179; b = 8'd53;  #10 
a = 8'd179; b = 8'd54;  #10 
a = 8'd179; b = 8'd55;  #10 
a = 8'd179; b = 8'd56;  #10 
a = 8'd179; b = 8'd57;  #10 
a = 8'd179; b = 8'd58;  #10 
a = 8'd179; b = 8'd59;  #10 
a = 8'd179; b = 8'd60;  #10 
a = 8'd179; b = 8'd61;  #10 
a = 8'd179; b = 8'd62;  #10 
a = 8'd179; b = 8'd63;  #10 
a = 8'd179; b = 8'd64;  #10 
a = 8'd179; b = 8'd65;  #10 
a = 8'd179; b = 8'd66;  #10 
a = 8'd179; b = 8'd67;  #10 
a = 8'd179; b = 8'd68;  #10 
a = 8'd179; b = 8'd69;  #10 
a = 8'd179; b = 8'd70;  #10 
a = 8'd179; b = 8'd71;  #10 
a = 8'd179; b = 8'd72;  #10 
a = 8'd179; b = 8'd73;  #10 
a = 8'd179; b = 8'd74;  #10 
a = 8'd179; b = 8'd75;  #10 
a = 8'd179; b = 8'd76;  #10 
a = 8'd179; b = 8'd77;  #10 
a = 8'd179; b = 8'd78;  #10 
a = 8'd179; b = 8'd79;  #10 
a = 8'd179; b = 8'd80;  #10 
a = 8'd179; b = 8'd81;  #10 
a = 8'd179; b = 8'd82;  #10 
a = 8'd179; b = 8'd83;  #10 
a = 8'd179; b = 8'd84;  #10 
a = 8'd179; b = 8'd85;  #10 
a = 8'd179; b = 8'd86;  #10 
a = 8'd179; b = 8'd87;  #10 
a = 8'd179; b = 8'd88;  #10 
a = 8'd179; b = 8'd89;  #10 
a = 8'd179; b = 8'd90;  #10 
a = 8'd179; b = 8'd91;  #10 
a = 8'd179; b = 8'd92;  #10 
a = 8'd179; b = 8'd93;  #10 
a = 8'd179; b = 8'd94;  #10 
a = 8'd179; b = 8'd95;  #10 
a = 8'd179; b = 8'd96;  #10 
a = 8'd179; b = 8'd97;  #10 
a = 8'd179; b = 8'd98;  #10 
a = 8'd179; b = 8'd99;  #10 
a = 8'd179; b = 8'd100;  #10 
a = 8'd179; b = 8'd101;  #10 
a = 8'd179; b = 8'd102;  #10 
a = 8'd179; b = 8'd103;  #10 
a = 8'd179; b = 8'd104;  #10 
a = 8'd179; b = 8'd105;  #10 
a = 8'd179; b = 8'd106;  #10 
a = 8'd179; b = 8'd107;  #10 
a = 8'd179; b = 8'd108;  #10 
a = 8'd179; b = 8'd109;  #10 
a = 8'd179; b = 8'd110;  #10 
a = 8'd179; b = 8'd111;  #10 
a = 8'd179; b = 8'd112;  #10 
a = 8'd179; b = 8'd113;  #10 
a = 8'd179; b = 8'd114;  #10 
a = 8'd179; b = 8'd115;  #10 
a = 8'd179; b = 8'd116;  #10 
a = 8'd179; b = 8'd117;  #10 
a = 8'd179; b = 8'd118;  #10 
a = 8'd179; b = 8'd119;  #10 
a = 8'd179; b = 8'd120;  #10 
a = 8'd179; b = 8'd121;  #10 
a = 8'd179; b = 8'd122;  #10 
a = 8'd179; b = 8'd123;  #10 
a = 8'd179; b = 8'd124;  #10 
a = 8'd179; b = 8'd125;  #10 
a = 8'd179; b = 8'd126;  #10 
a = 8'd179; b = 8'd127;  #10 
a = 8'd179; b = 8'd128;  #10 
a = 8'd179; b = 8'd129;  #10 
a = 8'd179; b = 8'd130;  #10 
a = 8'd179; b = 8'd131;  #10 
a = 8'd179; b = 8'd132;  #10 
a = 8'd179; b = 8'd133;  #10 
a = 8'd179; b = 8'd134;  #10 
a = 8'd179; b = 8'd135;  #10 
a = 8'd179; b = 8'd136;  #10 
a = 8'd179; b = 8'd137;  #10 
a = 8'd179; b = 8'd138;  #10 
a = 8'd179; b = 8'd139;  #10 
a = 8'd179; b = 8'd140;  #10 
a = 8'd179; b = 8'd141;  #10 
a = 8'd179; b = 8'd142;  #10 
a = 8'd179; b = 8'd143;  #10 
a = 8'd179; b = 8'd144;  #10 
a = 8'd179; b = 8'd145;  #10 
a = 8'd179; b = 8'd146;  #10 
a = 8'd179; b = 8'd147;  #10 
a = 8'd179; b = 8'd148;  #10 
a = 8'd179; b = 8'd149;  #10 
a = 8'd179; b = 8'd150;  #10 
a = 8'd179; b = 8'd151;  #10 
a = 8'd179; b = 8'd152;  #10 
a = 8'd179; b = 8'd153;  #10 
a = 8'd179; b = 8'd154;  #10 
a = 8'd179; b = 8'd155;  #10 
a = 8'd179; b = 8'd156;  #10 
a = 8'd179; b = 8'd157;  #10 
a = 8'd179; b = 8'd158;  #10 
a = 8'd179; b = 8'd159;  #10 
a = 8'd179; b = 8'd160;  #10 
a = 8'd179; b = 8'd161;  #10 
a = 8'd179; b = 8'd162;  #10 
a = 8'd179; b = 8'd163;  #10 
a = 8'd179; b = 8'd164;  #10 
a = 8'd179; b = 8'd165;  #10 
a = 8'd179; b = 8'd166;  #10 
a = 8'd179; b = 8'd167;  #10 
a = 8'd179; b = 8'd168;  #10 
a = 8'd179; b = 8'd169;  #10 
a = 8'd179; b = 8'd170;  #10 
a = 8'd179; b = 8'd171;  #10 
a = 8'd179; b = 8'd172;  #10 
a = 8'd179; b = 8'd173;  #10 
a = 8'd179; b = 8'd174;  #10 
a = 8'd179; b = 8'd175;  #10 
a = 8'd179; b = 8'd176;  #10 
a = 8'd179; b = 8'd177;  #10 
a = 8'd179; b = 8'd178;  #10 
a = 8'd179; b = 8'd179;  #10 
a = 8'd179; b = 8'd180;  #10 
a = 8'd179; b = 8'd181;  #10 
a = 8'd179; b = 8'd182;  #10 
a = 8'd179; b = 8'd183;  #10 
a = 8'd179; b = 8'd184;  #10 
a = 8'd179; b = 8'd185;  #10 
a = 8'd179; b = 8'd186;  #10 
a = 8'd179; b = 8'd187;  #10 
a = 8'd179; b = 8'd188;  #10 
a = 8'd179; b = 8'd189;  #10 
a = 8'd179; b = 8'd190;  #10 
a = 8'd179; b = 8'd191;  #10 
a = 8'd179; b = 8'd192;  #10 
a = 8'd179; b = 8'd193;  #10 
a = 8'd179; b = 8'd194;  #10 
a = 8'd179; b = 8'd195;  #10 
a = 8'd179; b = 8'd196;  #10 
a = 8'd179; b = 8'd197;  #10 
a = 8'd179; b = 8'd198;  #10 
a = 8'd179; b = 8'd199;  #10 
a = 8'd179; b = 8'd200;  #10 
a = 8'd179; b = 8'd201;  #10 
a = 8'd179; b = 8'd202;  #10 
a = 8'd179; b = 8'd203;  #10 
a = 8'd179; b = 8'd204;  #10 
a = 8'd179; b = 8'd205;  #10 
a = 8'd179; b = 8'd206;  #10 
a = 8'd179; b = 8'd207;  #10 
a = 8'd179; b = 8'd208;  #10 
a = 8'd179; b = 8'd209;  #10 
a = 8'd179; b = 8'd210;  #10 
a = 8'd179; b = 8'd211;  #10 
a = 8'd179; b = 8'd212;  #10 
a = 8'd179; b = 8'd213;  #10 
a = 8'd179; b = 8'd214;  #10 
a = 8'd179; b = 8'd215;  #10 
a = 8'd179; b = 8'd216;  #10 
a = 8'd179; b = 8'd217;  #10 
a = 8'd179; b = 8'd218;  #10 
a = 8'd179; b = 8'd219;  #10 
a = 8'd179; b = 8'd220;  #10 
a = 8'd179; b = 8'd221;  #10 
a = 8'd179; b = 8'd222;  #10 
a = 8'd179; b = 8'd223;  #10 
a = 8'd179; b = 8'd224;  #10 
a = 8'd179; b = 8'd225;  #10 
a = 8'd179; b = 8'd226;  #10 
a = 8'd179; b = 8'd227;  #10 
a = 8'd179; b = 8'd228;  #10 
a = 8'd179; b = 8'd229;  #10 
a = 8'd179; b = 8'd230;  #10 
a = 8'd179; b = 8'd231;  #10 
a = 8'd179; b = 8'd232;  #10 
a = 8'd179; b = 8'd233;  #10 
a = 8'd179; b = 8'd234;  #10 
a = 8'd179; b = 8'd235;  #10 
a = 8'd179; b = 8'd236;  #10 
a = 8'd179; b = 8'd237;  #10 
a = 8'd179; b = 8'd238;  #10 
a = 8'd179; b = 8'd239;  #10 
a = 8'd179; b = 8'd240;  #10 
a = 8'd179; b = 8'd241;  #10 
a = 8'd179; b = 8'd242;  #10 
a = 8'd179; b = 8'd243;  #10 
a = 8'd179; b = 8'd244;  #10 
a = 8'd179; b = 8'd245;  #10 
a = 8'd179; b = 8'd246;  #10 
a = 8'd179; b = 8'd247;  #10 
a = 8'd179; b = 8'd248;  #10 
a = 8'd179; b = 8'd249;  #10 
a = 8'd179; b = 8'd250;  #10 
a = 8'd179; b = 8'd251;  #10 
a = 8'd179; b = 8'd252;  #10 
a = 8'd179; b = 8'd253;  #10 
a = 8'd179; b = 8'd254;  #10 
a = 8'd179; b = 8'd255;  #10 
a = 8'd180; b = 8'd0;  #10 
a = 8'd180; b = 8'd1;  #10 
a = 8'd180; b = 8'd2;  #10 
a = 8'd180; b = 8'd3;  #10 
a = 8'd180; b = 8'd4;  #10 
a = 8'd180; b = 8'd5;  #10 
a = 8'd180; b = 8'd6;  #10 
a = 8'd180; b = 8'd7;  #10 
a = 8'd180; b = 8'd8;  #10 
a = 8'd180; b = 8'd9;  #10 
a = 8'd180; b = 8'd10;  #10 
a = 8'd180; b = 8'd11;  #10 
a = 8'd180; b = 8'd12;  #10 
a = 8'd180; b = 8'd13;  #10 
a = 8'd180; b = 8'd14;  #10 
a = 8'd180; b = 8'd15;  #10 
a = 8'd180; b = 8'd16;  #10 
a = 8'd180; b = 8'd17;  #10 
a = 8'd180; b = 8'd18;  #10 
a = 8'd180; b = 8'd19;  #10 
a = 8'd180; b = 8'd20;  #10 
a = 8'd180; b = 8'd21;  #10 
a = 8'd180; b = 8'd22;  #10 
a = 8'd180; b = 8'd23;  #10 
a = 8'd180; b = 8'd24;  #10 
a = 8'd180; b = 8'd25;  #10 
a = 8'd180; b = 8'd26;  #10 
a = 8'd180; b = 8'd27;  #10 
a = 8'd180; b = 8'd28;  #10 
a = 8'd180; b = 8'd29;  #10 
a = 8'd180; b = 8'd30;  #10 
a = 8'd180; b = 8'd31;  #10 
a = 8'd180; b = 8'd32;  #10 
a = 8'd180; b = 8'd33;  #10 
a = 8'd180; b = 8'd34;  #10 
a = 8'd180; b = 8'd35;  #10 
a = 8'd180; b = 8'd36;  #10 
a = 8'd180; b = 8'd37;  #10 
a = 8'd180; b = 8'd38;  #10 
a = 8'd180; b = 8'd39;  #10 
a = 8'd180; b = 8'd40;  #10 
a = 8'd180; b = 8'd41;  #10 
a = 8'd180; b = 8'd42;  #10 
a = 8'd180; b = 8'd43;  #10 
a = 8'd180; b = 8'd44;  #10 
a = 8'd180; b = 8'd45;  #10 
a = 8'd180; b = 8'd46;  #10 
a = 8'd180; b = 8'd47;  #10 
a = 8'd180; b = 8'd48;  #10 
a = 8'd180; b = 8'd49;  #10 
a = 8'd180; b = 8'd50;  #10 
a = 8'd180; b = 8'd51;  #10 
a = 8'd180; b = 8'd52;  #10 
a = 8'd180; b = 8'd53;  #10 
a = 8'd180; b = 8'd54;  #10 
a = 8'd180; b = 8'd55;  #10 
a = 8'd180; b = 8'd56;  #10 
a = 8'd180; b = 8'd57;  #10 
a = 8'd180; b = 8'd58;  #10 
a = 8'd180; b = 8'd59;  #10 
a = 8'd180; b = 8'd60;  #10 
a = 8'd180; b = 8'd61;  #10 
a = 8'd180; b = 8'd62;  #10 
a = 8'd180; b = 8'd63;  #10 
a = 8'd180; b = 8'd64;  #10 
a = 8'd180; b = 8'd65;  #10 
a = 8'd180; b = 8'd66;  #10 
a = 8'd180; b = 8'd67;  #10 
a = 8'd180; b = 8'd68;  #10 
a = 8'd180; b = 8'd69;  #10 
a = 8'd180; b = 8'd70;  #10 
a = 8'd180; b = 8'd71;  #10 
a = 8'd180; b = 8'd72;  #10 
a = 8'd180; b = 8'd73;  #10 
a = 8'd180; b = 8'd74;  #10 
a = 8'd180; b = 8'd75;  #10 
a = 8'd180; b = 8'd76;  #10 
a = 8'd180; b = 8'd77;  #10 
a = 8'd180; b = 8'd78;  #10 
a = 8'd180; b = 8'd79;  #10 
a = 8'd180; b = 8'd80;  #10 
a = 8'd180; b = 8'd81;  #10 
a = 8'd180; b = 8'd82;  #10 
a = 8'd180; b = 8'd83;  #10 
a = 8'd180; b = 8'd84;  #10 
a = 8'd180; b = 8'd85;  #10 
a = 8'd180; b = 8'd86;  #10 
a = 8'd180; b = 8'd87;  #10 
a = 8'd180; b = 8'd88;  #10 
a = 8'd180; b = 8'd89;  #10 
a = 8'd180; b = 8'd90;  #10 
a = 8'd180; b = 8'd91;  #10 
a = 8'd180; b = 8'd92;  #10 
a = 8'd180; b = 8'd93;  #10 
a = 8'd180; b = 8'd94;  #10 
a = 8'd180; b = 8'd95;  #10 
a = 8'd180; b = 8'd96;  #10 
a = 8'd180; b = 8'd97;  #10 
a = 8'd180; b = 8'd98;  #10 
a = 8'd180; b = 8'd99;  #10 
a = 8'd180; b = 8'd100;  #10 
a = 8'd180; b = 8'd101;  #10 
a = 8'd180; b = 8'd102;  #10 
a = 8'd180; b = 8'd103;  #10 
a = 8'd180; b = 8'd104;  #10 
a = 8'd180; b = 8'd105;  #10 
a = 8'd180; b = 8'd106;  #10 
a = 8'd180; b = 8'd107;  #10 
a = 8'd180; b = 8'd108;  #10 
a = 8'd180; b = 8'd109;  #10 
a = 8'd180; b = 8'd110;  #10 
a = 8'd180; b = 8'd111;  #10 
a = 8'd180; b = 8'd112;  #10 
a = 8'd180; b = 8'd113;  #10 
a = 8'd180; b = 8'd114;  #10 
a = 8'd180; b = 8'd115;  #10 
a = 8'd180; b = 8'd116;  #10 
a = 8'd180; b = 8'd117;  #10 
a = 8'd180; b = 8'd118;  #10 
a = 8'd180; b = 8'd119;  #10 
a = 8'd180; b = 8'd120;  #10 
a = 8'd180; b = 8'd121;  #10 
a = 8'd180; b = 8'd122;  #10 
a = 8'd180; b = 8'd123;  #10 
a = 8'd180; b = 8'd124;  #10 
a = 8'd180; b = 8'd125;  #10 
a = 8'd180; b = 8'd126;  #10 
a = 8'd180; b = 8'd127;  #10 
a = 8'd180; b = 8'd128;  #10 
a = 8'd180; b = 8'd129;  #10 
a = 8'd180; b = 8'd130;  #10 
a = 8'd180; b = 8'd131;  #10 
a = 8'd180; b = 8'd132;  #10 
a = 8'd180; b = 8'd133;  #10 
a = 8'd180; b = 8'd134;  #10 
a = 8'd180; b = 8'd135;  #10 
a = 8'd180; b = 8'd136;  #10 
a = 8'd180; b = 8'd137;  #10 
a = 8'd180; b = 8'd138;  #10 
a = 8'd180; b = 8'd139;  #10 
a = 8'd180; b = 8'd140;  #10 
a = 8'd180; b = 8'd141;  #10 
a = 8'd180; b = 8'd142;  #10 
a = 8'd180; b = 8'd143;  #10 
a = 8'd180; b = 8'd144;  #10 
a = 8'd180; b = 8'd145;  #10 
a = 8'd180; b = 8'd146;  #10 
a = 8'd180; b = 8'd147;  #10 
a = 8'd180; b = 8'd148;  #10 
a = 8'd180; b = 8'd149;  #10 
a = 8'd180; b = 8'd150;  #10 
a = 8'd180; b = 8'd151;  #10 
a = 8'd180; b = 8'd152;  #10 
a = 8'd180; b = 8'd153;  #10 
a = 8'd180; b = 8'd154;  #10 
a = 8'd180; b = 8'd155;  #10 
a = 8'd180; b = 8'd156;  #10 
a = 8'd180; b = 8'd157;  #10 
a = 8'd180; b = 8'd158;  #10 
a = 8'd180; b = 8'd159;  #10 
a = 8'd180; b = 8'd160;  #10 
a = 8'd180; b = 8'd161;  #10 
a = 8'd180; b = 8'd162;  #10 
a = 8'd180; b = 8'd163;  #10 
a = 8'd180; b = 8'd164;  #10 
a = 8'd180; b = 8'd165;  #10 
a = 8'd180; b = 8'd166;  #10 
a = 8'd180; b = 8'd167;  #10 
a = 8'd180; b = 8'd168;  #10 
a = 8'd180; b = 8'd169;  #10 
a = 8'd180; b = 8'd170;  #10 
a = 8'd180; b = 8'd171;  #10 
a = 8'd180; b = 8'd172;  #10 
a = 8'd180; b = 8'd173;  #10 
a = 8'd180; b = 8'd174;  #10 
a = 8'd180; b = 8'd175;  #10 
a = 8'd180; b = 8'd176;  #10 
a = 8'd180; b = 8'd177;  #10 
a = 8'd180; b = 8'd178;  #10 
a = 8'd180; b = 8'd179;  #10 
a = 8'd180; b = 8'd180;  #10 
a = 8'd180; b = 8'd181;  #10 
a = 8'd180; b = 8'd182;  #10 
a = 8'd180; b = 8'd183;  #10 
a = 8'd180; b = 8'd184;  #10 
a = 8'd180; b = 8'd185;  #10 
a = 8'd180; b = 8'd186;  #10 
a = 8'd180; b = 8'd187;  #10 
a = 8'd180; b = 8'd188;  #10 
a = 8'd180; b = 8'd189;  #10 
a = 8'd180; b = 8'd190;  #10 
a = 8'd180; b = 8'd191;  #10 
a = 8'd180; b = 8'd192;  #10 
a = 8'd180; b = 8'd193;  #10 
a = 8'd180; b = 8'd194;  #10 
a = 8'd180; b = 8'd195;  #10 
a = 8'd180; b = 8'd196;  #10 
a = 8'd180; b = 8'd197;  #10 
a = 8'd180; b = 8'd198;  #10 
a = 8'd180; b = 8'd199;  #10 
a = 8'd180; b = 8'd200;  #10 
a = 8'd180; b = 8'd201;  #10 
a = 8'd180; b = 8'd202;  #10 
a = 8'd180; b = 8'd203;  #10 
a = 8'd180; b = 8'd204;  #10 
a = 8'd180; b = 8'd205;  #10 
a = 8'd180; b = 8'd206;  #10 
a = 8'd180; b = 8'd207;  #10 
a = 8'd180; b = 8'd208;  #10 
a = 8'd180; b = 8'd209;  #10 
a = 8'd180; b = 8'd210;  #10 
a = 8'd180; b = 8'd211;  #10 
a = 8'd180; b = 8'd212;  #10 
a = 8'd180; b = 8'd213;  #10 
a = 8'd180; b = 8'd214;  #10 
a = 8'd180; b = 8'd215;  #10 
a = 8'd180; b = 8'd216;  #10 
a = 8'd180; b = 8'd217;  #10 
a = 8'd180; b = 8'd218;  #10 
a = 8'd180; b = 8'd219;  #10 
a = 8'd180; b = 8'd220;  #10 
a = 8'd180; b = 8'd221;  #10 
a = 8'd180; b = 8'd222;  #10 
a = 8'd180; b = 8'd223;  #10 
a = 8'd180; b = 8'd224;  #10 
a = 8'd180; b = 8'd225;  #10 
a = 8'd180; b = 8'd226;  #10 
a = 8'd180; b = 8'd227;  #10 
a = 8'd180; b = 8'd228;  #10 
a = 8'd180; b = 8'd229;  #10 
a = 8'd180; b = 8'd230;  #10 
a = 8'd180; b = 8'd231;  #10 
a = 8'd180; b = 8'd232;  #10 
a = 8'd180; b = 8'd233;  #10 
a = 8'd180; b = 8'd234;  #10 
a = 8'd180; b = 8'd235;  #10 
a = 8'd180; b = 8'd236;  #10 
a = 8'd180; b = 8'd237;  #10 
a = 8'd180; b = 8'd238;  #10 
a = 8'd180; b = 8'd239;  #10 
a = 8'd180; b = 8'd240;  #10 
a = 8'd180; b = 8'd241;  #10 
a = 8'd180; b = 8'd242;  #10 
a = 8'd180; b = 8'd243;  #10 
a = 8'd180; b = 8'd244;  #10 
a = 8'd180; b = 8'd245;  #10 
a = 8'd180; b = 8'd246;  #10 
a = 8'd180; b = 8'd247;  #10 
a = 8'd180; b = 8'd248;  #10 
a = 8'd180; b = 8'd249;  #10 
a = 8'd180; b = 8'd250;  #10 
a = 8'd180; b = 8'd251;  #10 
a = 8'd180; b = 8'd252;  #10 
a = 8'd180; b = 8'd253;  #10 
a = 8'd180; b = 8'd254;  #10 
a = 8'd180; b = 8'd255;  #10 
a = 8'd181; b = 8'd0;  #10 
a = 8'd181; b = 8'd1;  #10 
a = 8'd181; b = 8'd2;  #10 
a = 8'd181; b = 8'd3;  #10 
a = 8'd181; b = 8'd4;  #10 
a = 8'd181; b = 8'd5;  #10 
a = 8'd181; b = 8'd6;  #10 
a = 8'd181; b = 8'd7;  #10 
a = 8'd181; b = 8'd8;  #10 
a = 8'd181; b = 8'd9;  #10 
a = 8'd181; b = 8'd10;  #10 
a = 8'd181; b = 8'd11;  #10 
a = 8'd181; b = 8'd12;  #10 
a = 8'd181; b = 8'd13;  #10 
a = 8'd181; b = 8'd14;  #10 
a = 8'd181; b = 8'd15;  #10 
a = 8'd181; b = 8'd16;  #10 
a = 8'd181; b = 8'd17;  #10 
a = 8'd181; b = 8'd18;  #10 
a = 8'd181; b = 8'd19;  #10 
a = 8'd181; b = 8'd20;  #10 
a = 8'd181; b = 8'd21;  #10 
a = 8'd181; b = 8'd22;  #10 
a = 8'd181; b = 8'd23;  #10 
a = 8'd181; b = 8'd24;  #10 
a = 8'd181; b = 8'd25;  #10 
a = 8'd181; b = 8'd26;  #10 
a = 8'd181; b = 8'd27;  #10 
a = 8'd181; b = 8'd28;  #10 
a = 8'd181; b = 8'd29;  #10 
a = 8'd181; b = 8'd30;  #10 
a = 8'd181; b = 8'd31;  #10 
a = 8'd181; b = 8'd32;  #10 
a = 8'd181; b = 8'd33;  #10 
a = 8'd181; b = 8'd34;  #10 
a = 8'd181; b = 8'd35;  #10 
a = 8'd181; b = 8'd36;  #10 
a = 8'd181; b = 8'd37;  #10 
a = 8'd181; b = 8'd38;  #10 
a = 8'd181; b = 8'd39;  #10 
a = 8'd181; b = 8'd40;  #10 
a = 8'd181; b = 8'd41;  #10 
a = 8'd181; b = 8'd42;  #10 
a = 8'd181; b = 8'd43;  #10 
a = 8'd181; b = 8'd44;  #10 
a = 8'd181; b = 8'd45;  #10 
a = 8'd181; b = 8'd46;  #10 
a = 8'd181; b = 8'd47;  #10 
a = 8'd181; b = 8'd48;  #10 
a = 8'd181; b = 8'd49;  #10 
a = 8'd181; b = 8'd50;  #10 
a = 8'd181; b = 8'd51;  #10 
a = 8'd181; b = 8'd52;  #10 
a = 8'd181; b = 8'd53;  #10 
a = 8'd181; b = 8'd54;  #10 
a = 8'd181; b = 8'd55;  #10 
a = 8'd181; b = 8'd56;  #10 
a = 8'd181; b = 8'd57;  #10 
a = 8'd181; b = 8'd58;  #10 
a = 8'd181; b = 8'd59;  #10 
a = 8'd181; b = 8'd60;  #10 
a = 8'd181; b = 8'd61;  #10 
a = 8'd181; b = 8'd62;  #10 
a = 8'd181; b = 8'd63;  #10 
a = 8'd181; b = 8'd64;  #10 
a = 8'd181; b = 8'd65;  #10 
a = 8'd181; b = 8'd66;  #10 
a = 8'd181; b = 8'd67;  #10 
a = 8'd181; b = 8'd68;  #10 
a = 8'd181; b = 8'd69;  #10 
a = 8'd181; b = 8'd70;  #10 
a = 8'd181; b = 8'd71;  #10 
a = 8'd181; b = 8'd72;  #10 
a = 8'd181; b = 8'd73;  #10 
a = 8'd181; b = 8'd74;  #10 
a = 8'd181; b = 8'd75;  #10 
a = 8'd181; b = 8'd76;  #10 
a = 8'd181; b = 8'd77;  #10 
a = 8'd181; b = 8'd78;  #10 
a = 8'd181; b = 8'd79;  #10 
a = 8'd181; b = 8'd80;  #10 
a = 8'd181; b = 8'd81;  #10 
a = 8'd181; b = 8'd82;  #10 
a = 8'd181; b = 8'd83;  #10 
a = 8'd181; b = 8'd84;  #10 
a = 8'd181; b = 8'd85;  #10 
a = 8'd181; b = 8'd86;  #10 
a = 8'd181; b = 8'd87;  #10 
a = 8'd181; b = 8'd88;  #10 
a = 8'd181; b = 8'd89;  #10 
a = 8'd181; b = 8'd90;  #10 
a = 8'd181; b = 8'd91;  #10 
a = 8'd181; b = 8'd92;  #10 
a = 8'd181; b = 8'd93;  #10 
a = 8'd181; b = 8'd94;  #10 
a = 8'd181; b = 8'd95;  #10 
a = 8'd181; b = 8'd96;  #10 
a = 8'd181; b = 8'd97;  #10 
a = 8'd181; b = 8'd98;  #10 
a = 8'd181; b = 8'd99;  #10 
a = 8'd181; b = 8'd100;  #10 
a = 8'd181; b = 8'd101;  #10 
a = 8'd181; b = 8'd102;  #10 
a = 8'd181; b = 8'd103;  #10 
a = 8'd181; b = 8'd104;  #10 
a = 8'd181; b = 8'd105;  #10 
a = 8'd181; b = 8'd106;  #10 
a = 8'd181; b = 8'd107;  #10 
a = 8'd181; b = 8'd108;  #10 
a = 8'd181; b = 8'd109;  #10 
a = 8'd181; b = 8'd110;  #10 
a = 8'd181; b = 8'd111;  #10 
a = 8'd181; b = 8'd112;  #10 
a = 8'd181; b = 8'd113;  #10 
a = 8'd181; b = 8'd114;  #10 
a = 8'd181; b = 8'd115;  #10 
a = 8'd181; b = 8'd116;  #10 
a = 8'd181; b = 8'd117;  #10 
a = 8'd181; b = 8'd118;  #10 
a = 8'd181; b = 8'd119;  #10 
a = 8'd181; b = 8'd120;  #10 
a = 8'd181; b = 8'd121;  #10 
a = 8'd181; b = 8'd122;  #10 
a = 8'd181; b = 8'd123;  #10 
a = 8'd181; b = 8'd124;  #10 
a = 8'd181; b = 8'd125;  #10 
a = 8'd181; b = 8'd126;  #10 
a = 8'd181; b = 8'd127;  #10 
a = 8'd181; b = 8'd128;  #10 
a = 8'd181; b = 8'd129;  #10 
a = 8'd181; b = 8'd130;  #10 
a = 8'd181; b = 8'd131;  #10 
a = 8'd181; b = 8'd132;  #10 
a = 8'd181; b = 8'd133;  #10 
a = 8'd181; b = 8'd134;  #10 
a = 8'd181; b = 8'd135;  #10 
a = 8'd181; b = 8'd136;  #10 
a = 8'd181; b = 8'd137;  #10 
a = 8'd181; b = 8'd138;  #10 
a = 8'd181; b = 8'd139;  #10 
a = 8'd181; b = 8'd140;  #10 
a = 8'd181; b = 8'd141;  #10 
a = 8'd181; b = 8'd142;  #10 
a = 8'd181; b = 8'd143;  #10 
a = 8'd181; b = 8'd144;  #10 
a = 8'd181; b = 8'd145;  #10 
a = 8'd181; b = 8'd146;  #10 
a = 8'd181; b = 8'd147;  #10 
a = 8'd181; b = 8'd148;  #10 
a = 8'd181; b = 8'd149;  #10 
a = 8'd181; b = 8'd150;  #10 
a = 8'd181; b = 8'd151;  #10 
a = 8'd181; b = 8'd152;  #10 
a = 8'd181; b = 8'd153;  #10 
a = 8'd181; b = 8'd154;  #10 
a = 8'd181; b = 8'd155;  #10 
a = 8'd181; b = 8'd156;  #10 
a = 8'd181; b = 8'd157;  #10 
a = 8'd181; b = 8'd158;  #10 
a = 8'd181; b = 8'd159;  #10 
a = 8'd181; b = 8'd160;  #10 
a = 8'd181; b = 8'd161;  #10 
a = 8'd181; b = 8'd162;  #10 
a = 8'd181; b = 8'd163;  #10 
a = 8'd181; b = 8'd164;  #10 
a = 8'd181; b = 8'd165;  #10 
a = 8'd181; b = 8'd166;  #10 
a = 8'd181; b = 8'd167;  #10 
a = 8'd181; b = 8'd168;  #10 
a = 8'd181; b = 8'd169;  #10 
a = 8'd181; b = 8'd170;  #10 
a = 8'd181; b = 8'd171;  #10 
a = 8'd181; b = 8'd172;  #10 
a = 8'd181; b = 8'd173;  #10 
a = 8'd181; b = 8'd174;  #10 
a = 8'd181; b = 8'd175;  #10 
a = 8'd181; b = 8'd176;  #10 
a = 8'd181; b = 8'd177;  #10 
a = 8'd181; b = 8'd178;  #10 
a = 8'd181; b = 8'd179;  #10 
a = 8'd181; b = 8'd180;  #10 
a = 8'd181; b = 8'd181;  #10 
a = 8'd181; b = 8'd182;  #10 
a = 8'd181; b = 8'd183;  #10 
a = 8'd181; b = 8'd184;  #10 
a = 8'd181; b = 8'd185;  #10 
a = 8'd181; b = 8'd186;  #10 
a = 8'd181; b = 8'd187;  #10 
a = 8'd181; b = 8'd188;  #10 
a = 8'd181; b = 8'd189;  #10 
a = 8'd181; b = 8'd190;  #10 
a = 8'd181; b = 8'd191;  #10 
a = 8'd181; b = 8'd192;  #10 
a = 8'd181; b = 8'd193;  #10 
a = 8'd181; b = 8'd194;  #10 
a = 8'd181; b = 8'd195;  #10 
a = 8'd181; b = 8'd196;  #10 
a = 8'd181; b = 8'd197;  #10 
a = 8'd181; b = 8'd198;  #10 
a = 8'd181; b = 8'd199;  #10 
a = 8'd181; b = 8'd200;  #10 
a = 8'd181; b = 8'd201;  #10 
a = 8'd181; b = 8'd202;  #10 
a = 8'd181; b = 8'd203;  #10 
a = 8'd181; b = 8'd204;  #10 
a = 8'd181; b = 8'd205;  #10 
a = 8'd181; b = 8'd206;  #10 
a = 8'd181; b = 8'd207;  #10 
a = 8'd181; b = 8'd208;  #10 
a = 8'd181; b = 8'd209;  #10 
a = 8'd181; b = 8'd210;  #10 
a = 8'd181; b = 8'd211;  #10 
a = 8'd181; b = 8'd212;  #10 
a = 8'd181; b = 8'd213;  #10 
a = 8'd181; b = 8'd214;  #10 
a = 8'd181; b = 8'd215;  #10 
a = 8'd181; b = 8'd216;  #10 
a = 8'd181; b = 8'd217;  #10 
a = 8'd181; b = 8'd218;  #10 
a = 8'd181; b = 8'd219;  #10 
a = 8'd181; b = 8'd220;  #10 
a = 8'd181; b = 8'd221;  #10 
a = 8'd181; b = 8'd222;  #10 
a = 8'd181; b = 8'd223;  #10 
a = 8'd181; b = 8'd224;  #10 
a = 8'd181; b = 8'd225;  #10 
a = 8'd181; b = 8'd226;  #10 
a = 8'd181; b = 8'd227;  #10 
a = 8'd181; b = 8'd228;  #10 
a = 8'd181; b = 8'd229;  #10 
a = 8'd181; b = 8'd230;  #10 
a = 8'd181; b = 8'd231;  #10 
a = 8'd181; b = 8'd232;  #10 
a = 8'd181; b = 8'd233;  #10 
a = 8'd181; b = 8'd234;  #10 
a = 8'd181; b = 8'd235;  #10 
a = 8'd181; b = 8'd236;  #10 
a = 8'd181; b = 8'd237;  #10 
a = 8'd181; b = 8'd238;  #10 
a = 8'd181; b = 8'd239;  #10 
a = 8'd181; b = 8'd240;  #10 
a = 8'd181; b = 8'd241;  #10 
a = 8'd181; b = 8'd242;  #10 
a = 8'd181; b = 8'd243;  #10 
a = 8'd181; b = 8'd244;  #10 
a = 8'd181; b = 8'd245;  #10 
a = 8'd181; b = 8'd246;  #10 
a = 8'd181; b = 8'd247;  #10 
a = 8'd181; b = 8'd248;  #10 
a = 8'd181; b = 8'd249;  #10 
a = 8'd181; b = 8'd250;  #10 
a = 8'd181; b = 8'd251;  #10 
a = 8'd181; b = 8'd252;  #10 
a = 8'd181; b = 8'd253;  #10 
a = 8'd181; b = 8'd254;  #10 
a = 8'd181; b = 8'd255;  #10 
a = 8'd182; b = 8'd0;  #10 
a = 8'd182; b = 8'd1;  #10 
a = 8'd182; b = 8'd2;  #10 
a = 8'd182; b = 8'd3;  #10 
a = 8'd182; b = 8'd4;  #10 
a = 8'd182; b = 8'd5;  #10 
a = 8'd182; b = 8'd6;  #10 
a = 8'd182; b = 8'd7;  #10 
a = 8'd182; b = 8'd8;  #10 
a = 8'd182; b = 8'd9;  #10 
a = 8'd182; b = 8'd10;  #10 
a = 8'd182; b = 8'd11;  #10 
a = 8'd182; b = 8'd12;  #10 
a = 8'd182; b = 8'd13;  #10 
a = 8'd182; b = 8'd14;  #10 
a = 8'd182; b = 8'd15;  #10 
a = 8'd182; b = 8'd16;  #10 
a = 8'd182; b = 8'd17;  #10 
a = 8'd182; b = 8'd18;  #10 
a = 8'd182; b = 8'd19;  #10 
a = 8'd182; b = 8'd20;  #10 
a = 8'd182; b = 8'd21;  #10 
a = 8'd182; b = 8'd22;  #10 
a = 8'd182; b = 8'd23;  #10 
a = 8'd182; b = 8'd24;  #10 
a = 8'd182; b = 8'd25;  #10 
a = 8'd182; b = 8'd26;  #10 
a = 8'd182; b = 8'd27;  #10 
a = 8'd182; b = 8'd28;  #10 
a = 8'd182; b = 8'd29;  #10 
a = 8'd182; b = 8'd30;  #10 
a = 8'd182; b = 8'd31;  #10 
a = 8'd182; b = 8'd32;  #10 
a = 8'd182; b = 8'd33;  #10 
a = 8'd182; b = 8'd34;  #10 
a = 8'd182; b = 8'd35;  #10 
a = 8'd182; b = 8'd36;  #10 
a = 8'd182; b = 8'd37;  #10 
a = 8'd182; b = 8'd38;  #10 
a = 8'd182; b = 8'd39;  #10 
a = 8'd182; b = 8'd40;  #10 
a = 8'd182; b = 8'd41;  #10 
a = 8'd182; b = 8'd42;  #10 
a = 8'd182; b = 8'd43;  #10 
a = 8'd182; b = 8'd44;  #10 
a = 8'd182; b = 8'd45;  #10 
a = 8'd182; b = 8'd46;  #10 
a = 8'd182; b = 8'd47;  #10 
a = 8'd182; b = 8'd48;  #10 
a = 8'd182; b = 8'd49;  #10 
a = 8'd182; b = 8'd50;  #10 
a = 8'd182; b = 8'd51;  #10 
a = 8'd182; b = 8'd52;  #10 
a = 8'd182; b = 8'd53;  #10 
a = 8'd182; b = 8'd54;  #10 
a = 8'd182; b = 8'd55;  #10 
a = 8'd182; b = 8'd56;  #10 
a = 8'd182; b = 8'd57;  #10 
a = 8'd182; b = 8'd58;  #10 
a = 8'd182; b = 8'd59;  #10 
a = 8'd182; b = 8'd60;  #10 
a = 8'd182; b = 8'd61;  #10 
a = 8'd182; b = 8'd62;  #10 
a = 8'd182; b = 8'd63;  #10 
a = 8'd182; b = 8'd64;  #10 
a = 8'd182; b = 8'd65;  #10 
a = 8'd182; b = 8'd66;  #10 
a = 8'd182; b = 8'd67;  #10 
a = 8'd182; b = 8'd68;  #10 
a = 8'd182; b = 8'd69;  #10 
a = 8'd182; b = 8'd70;  #10 
a = 8'd182; b = 8'd71;  #10 
a = 8'd182; b = 8'd72;  #10 
a = 8'd182; b = 8'd73;  #10 
a = 8'd182; b = 8'd74;  #10 
a = 8'd182; b = 8'd75;  #10 
a = 8'd182; b = 8'd76;  #10 
a = 8'd182; b = 8'd77;  #10 
a = 8'd182; b = 8'd78;  #10 
a = 8'd182; b = 8'd79;  #10 
a = 8'd182; b = 8'd80;  #10 
a = 8'd182; b = 8'd81;  #10 
a = 8'd182; b = 8'd82;  #10 
a = 8'd182; b = 8'd83;  #10 
a = 8'd182; b = 8'd84;  #10 
a = 8'd182; b = 8'd85;  #10 
a = 8'd182; b = 8'd86;  #10 
a = 8'd182; b = 8'd87;  #10 
a = 8'd182; b = 8'd88;  #10 
a = 8'd182; b = 8'd89;  #10 
a = 8'd182; b = 8'd90;  #10 
a = 8'd182; b = 8'd91;  #10 
a = 8'd182; b = 8'd92;  #10 
a = 8'd182; b = 8'd93;  #10 
a = 8'd182; b = 8'd94;  #10 
a = 8'd182; b = 8'd95;  #10 
a = 8'd182; b = 8'd96;  #10 
a = 8'd182; b = 8'd97;  #10 
a = 8'd182; b = 8'd98;  #10 
a = 8'd182; b = 8'd99;  #10 
a = 8'd182; b = 8'd100;  #10 
a = 8'd182; b = 8'd101;  #10 
a = 8'd182; b = 8'd102;  #10 
a = 8'd182; b = 8'd103;  #10 
a = 8'd182; b = 8'd104;  #10 
a = 8'd182; b = 8'd105;  #10 
a = 8'd182; b = 8'd106;  #10 
a = 8'd182; b = 8'd107;  #10 
a = 8'd182; b = 8'd108;  #10 
a = 8'd182; b = 8'd109;  #10 
a = 8'd182; b = 8'd110;  #10 
a = 8'd182; b = 8'd111;  #10 
a = 8'd182; b = 8'd112;  #10 
a = 8'd182; b = 8'd113;  #10 
a = 8'd182; b = 8'd114;  #10 
a = 8'd182; b = 8'd115;  #10 
a = 8'd182; b = 8'd116;  #10 
a = 8'd182; b = 8'd117;  #10 
a = 8'd182; b = 8'd118;  #10 
a = 8'd182; b = 8'd119;  #10 
a = 8'd182; b = 8'd120;  #10 
a = 8'd182; b = 8'd121;  #10 
a = 8'd182; b = 8'd122;  #10 
a = 8'd182; b = 8'd123;  #10 
a = 8'd182; b = 8'd124;  #10 
a = 8'd182; b = 8'd125;  #10 
a = 8'd182; b = 8'd126;  #10 
a = 8'd182; b = 8'd127;  #10 
a = 8'd182; b = 8'd128;  #10 
a = 8'd182; b = 8'd129;  #10 
a = 8'd182; b = 8'd130;  #10 
a = 8'd182; b = 8'd131;  #10 
a = 8'd182; b = 8'd132;  #10 
a = 8'd182; b = 8'd133;  #10 
a = 8'd182; b = 8'd134;  #10 
a = 8'd182; b = 8'd135;  #10 
a = 8'd182; b = 8'd136;  #10 
a = 8'd182; b = 8'd137;  #10 
a = 8'd182; b = 8'd138;  #10 
a = 8'd182; b = 8'd139;  #10 
a = 8'd182; b = 8'd140;  #10 
a = 8'd182; b = 8'd141;  #10 
a = 8'd182; b = 8'd142;  #10 
a = 8'd182; b = 8'd143;  #10 
a = 8'd182; b = 8'd144;  #10 
a = 8'd182; b = 8'd145;  #10 
a = 8'd182; b = 8'd146;  #10 
a = 8'd182; b = 8'd147;  #10 
a = 8'd182; b = 8'd148;  #10 
a = 8'd182; b = 8'd149;  #10 
a = 8'd182; b = 8'd150;  #10 
a = 8'd182; b = 8'd151;  #10 
a = 8'd182; b = 8'd152;  #10 
a = 8'd182; b = 8'd153;  #10 
a = 8'd182; b = 8'd154;  #10 
a = 8'd182; b = 8'd155;  #10 
a = 8'd182; b = 8'd156;  #10 
a = 8'd182; b = 8'd157;  #10 
a = 8'd182; b = 8'd158;  #10 
a = 8'd182; b = 8'd159;  #10 
a = 8'd182; b = 8'd160;  #10 
a = 8'd182; b = 8'd161;  #10 
a = 8'd182; b = 8'd162;  #10 
a = 8'd182; b = 8'd163;  #10 
a = 8'd182; b = 8'd164;  #10 
a = 8'd182; b = 8'd165;  #10 
a = 8'd182; b = 8'd166;  #10 
a = 8'd182; b = 8'd167;  #10 
a = 8'd182; b = 8'd168;  #10 
a = 8'd182; b = 8'd169;  #10 
a = 8'd182; b = 8'd170;  #10 
a = 8'd182; b = 8'd171;  #10 
a = 8'd182; b = 8'd172;  #10 
a = 8'd182; b = 8'd173;  #10 
a = 8'd182; b = 8'd174;  #10 
a = 8'd182; b = 8'd175;  #10 
a = 8'd182; b = 8'd176;  #10 
a = 8'd182; b = 8'd177;  #10 
a = 8'd182; b = 8'd178;  #10 
a = 8'd182; b = 8'd179;  #10 
a = 8'd182; b = 8'd180;  #10 
a = 8'd182; b = 8'd181;  #10 
a = 8'd182; b = 8'd182;  #10 
a = 8'd182; b = 8'd183;  #10 
a = 8'd182; b = 8'd184;  #10 
a = 8'd182; b = 8'd185;  #10 
a = 8'd182; b = 8'd186;  #10 
a = 8'd182; b = 8'd187;  #10 
a = 8'd182; b = 8'd188;  #10 
a = 8'd182; b = 8'd189;  #10 
a = 8'd182; b = 8'd190;  #10 
a = 8'd182; b = 8'd191;  #10 
a = 8'd182; b = 8'd192;  #10 
a = 8'd182; b = 8'd193;  #10 
a = 8'd182; b = 8'd194;  #10 
a = 8'd182; b = 8'd195;  #10 
a = 8'd182; b = 8'd196;  #10 
a = 8'd182; b = 8'd197;  #10 
a = 8'd182; b = 8'd198;  #10 
a = 8'd182; b = 8'd199;  #10 
a = 8'd182; b = 8'd200;  #10 
a = 8'd182; b = 8'd201;  #10 
a = 8'd182; b = 8'd202;  #10 
a = 8'd182; b = 8'd203;  #10 
a = 8'd182; b = 8'd204;  #10 
a = 8'd182; b = 8'd205;  #10 
a = 8'd182; b = 8'd206;  #10 
a = 8'd182; b = 8'd207;  #10 
a = 8'd182; b = 8'd208;  #10 
a = 8'd182; b = 8'd209;  #10 
a = 8'd182; b = 8'd210;  #10 
a = 8'd182; b = 8'd211;  #10 
a = 8'd182; b = 8'd212;  #10 
a = 8'd182; b = 8'd213;  #10 
a = 8'd182; b = 8'd214;  #10 
a = 8'd182; b = 8'd215;  #10 
a = 8'd182; b = 8'd216;  #10 
a = 8'd182; b = 8'd217;  #10 
a = 8'd182; b = 8'd218;  #10 
a = 8'd182; b = 8'd219;  #10 
a = 8'd182; b = 8'd220;  #10 
a = 8'd182; b = 8'd221;  #10 
a = 8'd182; b = 8'd222;  #10 
a = 8'd182; b = 8'd223;  #10 
a = 8'd182; b = 8'd224;  #10 
a = 8'd182; b = 8'd225;  #10 
a = 8'd182; b = 8'd226;  #10 
a = 8'd182; b = 8'd227;  #10 
a = 8'd182; b = 8'd228;  #10 
a = 8'd182; b = 8'd229;  #10 
a = 8'd182; b = 8'd230;  #10 
a = 8'd182; b = 8'd231;  #10 
a = 8'd182; b = 8'd232;  #10 
a = 8'd182; b = 8'd233;  #10 
a = 8'd182; b = 8'd234;  #10 
a = 8'd182; b = 8'd235;  #10 
a = 8'd182; b = 8'd236;  #10 
a = 8'd182; b = 8'd237;  #10 
a = 8'd182; b = 8'd238;  #10 
a = 8'd182; b = 8'd239;  #10 
a = 8'd182; b = 8'd240;  #10 
a = 8'd182; b = 8'd241;  #10 
a = 8'd182; b = 8'd242;  #10 
a = 8'd182; b = 8'd243;  #10 
a = 8'd182; b = 8'd244;  #10 
a = 8'd182; b = 8'd245;  #10 
a = 8'd182; b = 8'd246;  #10 
a = 8'd182; b = 8'd247;  #10 
a = 8'd182; b = 8'd248;  #10 
a = 8'd182; b = 8'd249;  #10 
a = 8'd182; b = 8'd250;  #10 
a = 8'd182; b = 8'd251;  #10 
a = 8'd182; b = 8'd252;  #10 
a = 8'd182; b = 8'd253;  #10 
a = 8'd182; b = 8'd254;  #10 
a = 8'd182; b = 8'd255;  #10 
a = 8'd183; b = 8'd0;  #10 
a = 8'd183; b = 8'd1;  #10 
a = 8'd183; b = 8'd2;  #10 
a = 8'd183; b = 8'd3;  #10 
a = 8'd183; b = 8'd4;  #10 
a = 8'd183; b = 8'd5;  #10 
a = 8'd183; b = 8'd6;  #10 
a = 8'd183; b = 8'd7;  #10 
a = 8'd183; b = 8'd8;  #10 
a = 8'd183; b = 8'd9;  #10 
a = 8'd183; b = 8'd10;  #10 
a = 8'd183; b = 8'd11;  #10 
a = 8'd183; b = 8'd12;  #10 
a = 8'd183; b = 8'd13;  #10 
a = 8'd183; b = 8'd14;  #10 
a = 8'd183; b = 8'd15;  #10 
a = 8'd183; b = 8'd16;  #10 
a = 8'd183; b = 8'd17;  #10 
a = 8'd183; b = 8'd18;  #10 
a = 8'd183; b = 8'd19;  #10 
a = 8'd183; b = 8'd20;  #10 
a = 8'd183; b = 8'd21;  #10 
a = 8'd183; b = 8'd22;  #10 
a = 8'd183; b = 8'd23;  #10 
a = 8'd183; b = 8'd24;  #10 
a = 8'd183; b = 8'd25;  #10 
a = 8'd183; b = 8'd26;  #10 
a = 8'd183; b = 8'd27;  #10 
a = 8'd183; b = 8'd28;  #10 
a = 8'd183; b = 8'd29;  #10 
a = 8'd183; b = 8'd30;  #10 
a = 8'd183; b = 8'd31;  #10 
a = 8'd183; b = 8'd32;  #10 
a = 8'd183; b = 8'd33;  #10 
a = 8'd183; b = 8'd34;  #10 
a = 8'd183; b = 8'd35;  #10 
a = 8'd183; b = 8'd36;  #10 
a = 8'd183; b = 8'd37;  #10 
a = 8'd183; b = 8'd38;  #10 
a = 8'd183; b = 8'd39;  #10 
a = 8'd183; b = 8'd40;  #10 
a = 8'd183; b = 8'd41;  #10 
a = 8'd183; b = 8'd42;  #10 
a = 8'd183; b = 8'd43;  #10 
a = 8'd183; b = 8'd44;  #10 
a = 8'd183; b = 8'd45;  #10 
a = 8'd183; b = 8'd46;  #10 
a = 8'd183; b = 8'd47;  #10 
a = 8'd183; b = 8'd48;  #10 
a = 8'd183; b = 8'd49;  #10 
a = 8'd183; b = 8'd50;  #10 
a = 8'd183; b = 8'd51;  #10 
a = 8'd183; b = 8'd52;  #10 
a = 8'd183; b = 8'd53;  #10 
a = 8'd183; b = 8'd54;  #10 
a = 8'd183; b = 8'd55;  #10 
a = 8'd183; b = 8'd56;  #10 
a = 8'd183; b = 8'd57;  #10 
a = 8'd183; b = 8'd58;  #10 
a = 8'd183; b = 8'd59;  #10 
a = 8'd183; b = 8'd60;  #10 
a = 8'd183; b = 8'd61;  #10 
a = 8'd183; b = 8'd62;  #10 
a = 8'd183; b = 8'd63;  #10 
a = 8'd183; b = 8'd64;  #10 
a = 8'd183; b = 8'd65;  #10 
a = 8'd183; b = 8'd66;  #10 
a = 8'd183; b = 8'd67;  #10 
a = 8'd183; b = 8'd68;  #10 
a = 8'd183; b = 8'd69;  #10 
a = 8'd183; b = 8'd70;  #10 
a = 8'd183; b = 8'd71;  #10 
a = 8'd183; b = 8'd72;  #10 
a = 8'd183; b = 8'd73;  #10 
a = 8'd183; b = 8'd74;  #10 
a = 8'd183; b = 8'd75;  #10 
a = 8'd183; b = 8'd76;  #10 
a = 8'd183; b = 8'd77;  #10 
a = 8'd183; b = 8'd78;  #10 
a = 8'd183; b = 8'd79;  #10 
a = 8'd183; b = 8'd80;  #10 
a = 8'd183; b = 8'd81;  #10 
a = 8'd183; b = 8'd82;  #10 
a = 8'd183; b = 8'd83;  #10 
a = 8'd183; b = 8'd84;  #10 
a = 8'd183; b = 8'd85;  #10 
a = 8'd183; b = 8'd86;  #10 
a = 8'd183; b = 8'd87;  #10 
a = 8'd183; b = 8'd88;  #10 
a = 8'd183; b = 8'd89;  #10 
a = 8'd183; b = 8'd90;  #10 
a = 8'd183; b = 8'd91;  #10 
a = 8'd183; b = 8'd92;  #10 
a = 8'd183; b = 8'd93;  #10 
a = 8'd183; b = 8'd94;  #10 
a = 8'd183; b = 8'd95;  #10 
a = 8'd183; b = 8'd96;  #10 
a = 8'd183; b = 8'd97;  #10 
a = 8'd183; b = 8'd98;  #10 
a = 8'd183; b = 8'd99;  #10 
a = 8'd183; b = 8'd100;  #10 
a = 8'd183; b = 8'd101;  #10 
a = 8'd183; b = 8'd102;  #10 
a = 8'd183; b = 8'd103;  #10 
a = 8'd183; b = 8'd104;  #10 
a = 8'd183; b = 8'd105;  #10 
a = 8'd183; b = 8'd106;  #10 
a = 8'd183; b = 8'd107;  #10 
a = 8'd183; b = 8'd108;  #10 
a = 8'd183; b = 8'd109;  #10 
a = 8'd183; b = 8'd110;  #10 
a = 8'd183; b = 8'd111;  #10 
a = 8'd183; b = 8'd112;  #10 
a = 8'd183; b = 8'd113;  #10 
a = 8'd183; b = 8'd114;  #10 
a = 8'd183; b = 8'd115;  #10 
a = 8'd183; b = 8'd116;  #10 
a = 8'd183; b = 8'd117;  #10 
a = 8'd183; b = 8'd118;  #10 
a = 8'd183; b = 8'd119;  #10 
a = 8'd183; b = 8'd120;  #10 
a = 8'd183; b = 8'd121;  #10 
a = 8'd183; b = 8'd122;  #10 
a = 8'd183; b = 8'd123;  #10 
a = 8'd183; b = 8'd124;  #10 
a = 8'd183; b = 8'd125;  #10 
a = 8'd183; b = 8'd126;  #10 
a = 8'd183; b = 8'd127;  #10 
a = 8'd183; b = 8'd128;  #10 
a = 8'd183; b = 8'd129;  #10 
a = 8'd183; b = 8'd130;  #10 
a = 8'd183; b = 8'd131;  #10 
a = 8'd183; b = 8'd132;  #10 
a = 8'd183; b = 8'd133;  #10 
a = 8'd183; b = 8'd134;  #10 
a = 8'd183; b = 8'd135;  #10 
a = 8'd183; b = 8'd136;  #10 
a = 8'd183; b = 8'd137;  #10 
a = 8'd183; b = 8'd138;  #10 
a = 8'd183; b = 8'd139;  #10 
a = 8'd183; b = 8'd140;  #10 
a = 8'd183; b = 8'd141;  #10 
a = 8'd183; b = 8'd142;  #10 
a = 8'd183; b = 8'd143;  #10 
a = 8'd183; b = 8'd144;  #10 
a = 8'd183; b = 8'd145;  #10 
a = 8'd183; b = 8'd146;  #10 
a = 8'd183; b = 8'd147;  #10 
a = 8'd183; b = 8'd148;  #10 
a = 8'd183; b = 8'd149;  #10 
a = 8'd183; b = 8'd150;  #10 
a = 8'd183; b = 8'd151;  #10 
a = 8'd183; b = 8'd152;  #10 
a = 8'd183; b = 8'd153;  #10 
a = 8'd183; b = 8'd154;  #10 
a = 8'd183; b = 8'd155;  #10 
a = 8'd183; b = 8'd156;  #10 
a = 8'd183; b = 8'd157;  #10 
a = 8'd183; b = 8'd158;  #10 
a = 8'd183; b = 8'd159;  #10 
a = 8'd183; b = 8'd160;  #10 
a = 8'd183; b = 8'd161;  #10 
a = 8'd183; b = 8'd162;  #10 
a = 8'd183; b = 8'd163;  #10 
a = 8'd183; b = 8'd164;  #10 
a = 8'd183; b = 8'd165;  #10 
a = 8'd183; b = 8'd166;  #10 
a = 8'd183; b = 8'd167;  #10 
a = 8'd183; b = 8'd168;  #10 
a = 8'd183; b = 8'd169;  #10 
a = 8'd183; b = 8'd170;  #10 
a = 8'd183; b = 8'd171;  #10 
a = 8'd183; b = 8'd172;  #10 
a = 8'd183; b = 8'd173;  #10 
a = 8'd183; b = 8'd174;  #10 
a = 8'd183; b = 8'd175;  #10 
a = 8'd183; b = 8'd176;  #10 
a = 8'd183; b = 8'd177;  #10 
a = 8'd183; b = 8'd178;  #10 
a = 8'd183; b = 8'd179;  #10 
a = 8'd183; b = 8'd180;  #10 
a = 8'd183; b = 8'd181;  #10 
a = 8'd183; b = 8'd182;  #10 
a = 8'd183; b = 8'd183;  #10 
a = 8'd183; b = 8'd184;  #10 
a = 8'd183; b = 8'd185;  #10 
a = 8'd183; b = 8'd186;  #10 
a = 8'd183; b = 8'd187;  #10 
a = 8'd183; b = 8'd188;  #10 
a = 8'd183; b = 8'd189;  #10 
a = 8'd183; b = 8'd190;  #10 
a = 8'd183; b = 8'd191;  #10 
a = 8'd183; b = 8'd192;  #10 
a = 8'd183; b = 8'd193;  #10 
a = 8'd183; b = 8'd194;  #10 
a = 8'd183; b = 8'd195;  #10 
a = 8'd183; b = 8'd196;  #10 
a = 8'd183; b = 8'd197;  #10 
a = 8'd183; b = 8'd198;  #10 
a = 8'd183; b = 8'd199;  #10 
a = 8'd183; b = 8'd200;  #10 
a = 8'd183; b = 8'd201;  #10 
a = 8'd183; b = 8'd202;  #10 
a = 8'd183; b = 8'd203;  #10 
a = 8'd183; b = 8'd204;  #10 
a = 8'd183; b = 8'd205;  #10 
a = 8'd183; b = 8'd206;  #10 
a = 8'd183; b = 8'd207;  #10 
a = 8'd183; b = 8'd208;  #10 
a = 8'd183; b = 8'd209;  #10 
a = 8'd183; b = 8'd210;  #10 
a = 8'd183; b = 8'd211;  #10 
a = 8'd183; b = 8'd212;  #10 
a = 8'd183; b = 8'd213;  #10 
a = 8'd183; b = 8'd214;  #10 
a = 8'd183; b = 8'd215;  #10 
a = 8'd183; b = 8'd216;  #10 
a = 8'd183; b = 8'd217;  #10 
a = 8'd183; b = 8'd218;  #10 
a = 8'd183; b = 8'd219;  #10 
a = 8'd183; b = 8'd220;  #10 
a = 8'd183; b = 8'd221;  #10 
a = 8'd183; b = 8'd222;  #10 
a = 8'd183; b = 8'd223;  #10 
a = 8'd183; b = 8'd224;  #10 
a = 8'd183; b = 8'd225;  #10 
a = 8'd183; b = 8'd226;  #10 
a = 8'd183; b = 8'd227;  #10 
a = 8'd183; b = 8'd228;  #10 
a = 8'd183; b = 8'd229;  #10 
a = 8'd183; b = 8'd230;  #10 
a = 8'd183; b = 8'd231;  #10 
a = 8'd183; b = 8'd232;  #10 
a = 8'd183; b = 8'd233;  #10 
a = 8'd183; b = 8'd234;  #10 
a = 8'd183; b = 8'd235;  #10 
a = 8'd183; b = 8'd236;  #10 
a = 8'd183; b = 8'd237;  #10 
a = 8'd183; b = 8'd238;  #10 
a = 8'd183; b = 8'd239;  #10 
a = 8'd183; b = 8'd240;  #10 
a = 8'd183; b = 8'd241;  #10 
a = 8'd183; b = 8'd242;  #10 
a = 8'd183; b = 8'd243;  #10 
a = 8'd183; b = 8'd244;  #10 
a = 8'd183; b = 8'd245;  #10 
a = 8'd183; b = 8'd246;  #10 
a = 8'd183; b = 8'd247;  #10 
a = 8'd183; b = 8'd248;  #10 
a = 8'd183; b = 8'd249;  #10 
a = 8'd183; b = 8'd250;  #10 
a = 8'd183; b = 8'd251;  #10 
a = 8'd183; b = 8'd252;  #10 
a = 8'd183; b = 8'd253;  #10 
a = 8'd183; b = 8'd254;  #10 
a = 8'd183; b = 8'd255;  #10 
a = 8'd184; b = 8'd0;  #10 
a = 8'd184; b = 8'd1;  #10 
a = 8'd184; b = 8'd2;  #10 
a = 8'd184; b = 8'd3;  #10 
a = 8'd184; b = 8'd4;  #10 
a = 8'd184; b = 8'd5;  #10 
a = 8'd184; b = 8'd6;  #10 
a = 8'd184; b = 8'd7;  #10 
a = 8'd184; b = 8'd8;  #10 
a = 8'd184; b = 8'd9;  #10 
a = 8'd184; b = 8'd10;  #10 
a = 8'd184; b = 8'd11;  #10 
a = 8'd184; b = 8'd12;  #10 
a = 8'd184; b = 8'd13;  #10 
a = 8'd184; b = 8'd14;  #10 
a = 8'd184; b = 8'd15;  #10 
a = 8'd184; b = 8'd16;  #10 
a = 8'd184; b = 8'd17;  #10 
a = 8'd184; b = 8'd18;  #10 
a = 8'd184; b = 8'd19;  #10 
a = 8'd184; b = 8'd20;  #10 
a = 8'd184; b = 8'd21;  #10 
a = 8'd184; b = 8'd22;  #10 
a = 8'd184; b = 8'd23;  #10 
a = 8'd184; b = 8'd24;  #10 
a = 8'd184; b = 8'd25;  #10 
a = 8'd184; b = 8'd26;  #10 
a = 8'd184; b = 8'd27;  #10 
a = 8'd184; b = 8'd28;  #10 
a = 8'd184; b = 8'd29;  #10 
a = 8'd184; b = 8'd30;  #10 
a = 8'd184; b = 8'd31;  #10 
a = 8'd184; b = 8'd32;  #10 
a = 8'd184; b = 8'd33;  #10 
a = 8'd184; b = 8'd34;  #10 
a = 8'd184; b = 8'd35;  #10 
a = 8'd184; b = 8'd36;  #10 
a = 8'd184; b = 8'd37;  #10 
a = 8'd184; b = 8'd38;  #10 
a = 8'd184; b = 8'd39;  #10 
a = 8'd184; b = 8'd40;  #10 
a = 8'd184; b = 8'd41;  #10 
a = 8'd184; b = 8'd42;  #10 
a = 8'd184; b = 8'd43;  #10 
a = 8'd184; b = 8'd44;  #10 
a = 8'd184; b = 8'd45;  #10 
a = 8'd184; b = 8'd46;  #10 
a = 8'd184; b = 8'd47;  #10 
a = 8'd184; b = 8'd48;  #10 
a = 8'd184; b = 8'd49;  #10 
a = 8'd184; b = 8'd50;  #10 
a = 8'd184; b = 8'd51;  #10 
a = 8'd184; b = 8'd52;  #10 
a = 8'd184; b = 8'd53;  #10 
a = 8'd184; b = 8'd54;  #10 
a = 8'd184; b = 8'd55;  #10 
a = 8'd184; b = 8'd56;  #10 
a = 8'd184; b = 8'd57;  #10 
a = 8'd184; b = 8'd58;  #10 
a = 8'd184; b = 8'd59;  #10 
a = 8'd184; b = 8'd60;  #10 
a = 8'd184; b = 8'd61;  #10 
a = 8'd184; b = 8'd62;  #10 
a = 8'd184; b = 8'd63;  #10 
a = 8'd184; b = 8'd64;  #10 
a = 8'd184; b = 8'd65;  #10 
a = 8'd184; b = 8'd66;  #10 
a = 8'd184; b = 8'd67;  #10 
a = 8'd184; b = 8'd68;  #10 
a = 8'd184; b = 8'd69;  #10 
a = 8'd184; b = 8'd70;  #10 
a = 8'd184; b = 8'd71;  #10 
a = 8'd184; b = 8'd72;  #10 
a = 8'd184; b = 8'd73;  #10 
a = 8'd184; b = 8'd74;  #10 
a = 8'd184; b = 8'd75;  #10 
a = 8'd184; b = 8'd76;  #10 
a = 8'd184; b = 8'd77;  #10 
a = 8'd184; b = 8'd78;  #10 
a = 8'd184; b = 8'd79;  #10 
a = 8'd184; b = 8'd80;  #10 
a = 8'd184; b = 8'd81;  #10 
a = 8'd184; b = 8'd82;  #10 
a = 8'd184; b = 8'd83;  #10 
a = 8'd184; b = 8'd84;  #10 
a = 8'd184; b = 8'd85;  #10 
a = 8'd184; b = 8'd86;  #10 
a = 8'd184; b = 8'd87;  #10 
a = 8'd184; b = 8'd88;  #10 
a = 8'd184; b = 8'd89;  #10 
a = 8'd184; b = 8'd90;  #10 
a = 8'd184; b = 8'd91;  #10 
a = 8'd184; b = 8'd92;  #10 
a = 8'd184; b = 8'd93;  #10 
a = 8'd184; b = 8'd94;  #10 
a = 8'd184; b = 8'd95;  #10 
a = 8'd184; b = 8'd96;  #10 
a = 8'd184; b = 8'd97;  #10 
a = 8'd184; b = 8'd98;  #10 
a = 8'd184; b = 8'd99;  #10 
a = 8'd184; b = 8'd100;  #10 
a = 8'd184; b = 8'd101;  #10 
a = 8'd184; b = 8'd102;  #10 
a = 8'd184; b = 8'd103;  #10 
a = 8'd184; b = 8'd104;  #10 
a = 8'd184; b = 8'd105;  #10 
a = 8'd184; b = 8'd106;  #10 
a = 8'd184; b = 8'd107;  #10 
a = 8'd184; b = 8'd108;  #10 
a = 8'd184; b = 8'd109;  #10 
a = 8'd184; b = 8'd110;  #10 
a = 8'd184; b = 8'd111;  #10 
a = 8'd184; b = 8'd112;  #10 
a = 8'd184; b = 8'd113;  #10 
a = 8'd184; b = 8'd114;  #10 
a = 8'd184; b = 8'd115;  #10 
a = 8'd184; b = 8'd116;  #10 
a = 8'd184; b = 8'd117;  #10 
a = 8'd184; b = 8'd118;  #10 
a = 8'd184; b = 8'd119;  #10 
a = 8'd184; b = 8'd120;  #10 
a = 8'd184; b = 8'd121;  #10 
a = 8'd184; b = 8'd122;  #10 
a = 8'd184; b = 8'd123;  #10 
a = 8'd184; b = 8'd124;  #10 
a = 8'd184; b = 8'd125;  #10 
a = 8'd184; b = 8'd126;  #10 
a = 8'd184; b = 8'd127;  #10 
a = 8'd184; b = 8'd128;  #10 
a = 8'd184; b = 8'd129;  #10 
a = 8'd184; b = 8'd130;  #10 
a = 8'd184; b = 8'd131;  #10 
a = 8'd184; b = 8'd132;  #10 
a = 8'd184; b = 8'd133;  #10 
a = 8'd184; b = 8'd134;  #10 
a = 8'd184; b = 8'd135;  #10 
a = 8'd184; b = 8'd136;  #10 
a = 8'd184; b = 8'd137;  #10 
a = 8'd184; b = 8'd138;  #10 
a = 8'd184; b = 8'd139;  #10 
a = 8'd184; b = 8'd140;  #10 
a = 8'd184; b = 8'd141;  #10 
a = 8'd184; b = 8'd142;  #10 
a = 8'd184; b = 8'd143;  #10 
a = 8'd184; b = 8'd144;  #10 
a = 8'd184; b = 8'd145;  #10 
a = 8'd184; b = 8'd146;  #10 
a = 8'd184; b = 8'd147;  #10 
a = 8'd184; b = 8'd148;  #10 
a = 8'd184; b = 8'd149;  #10 
a = 8'd184; b = 8'd150;  #10 
a = 8'd184; b = 8'd151;  #10 
a = 8'd184; b = 8'd152;  #10 
a = 8'd184; b = 8'd153;  #10 
a = 8'd184; b = 8'd154;  #10 
a = 8'd184; b = 8'd155;  #10 
a = 8'd184; b = 8'd156;  #10 
a = 8'd184; b = 8'd157;  #10 
a = 8'd184; b = 8'd158;  #10 
a = 8'd184; b = 8'd159;  #10 
a = 8'd184; b = 8'd160;  #10 
a = 8'd184; b = 8'd161;  #10 
a = 8'd184; b = 8'd162;  #10 
a = 8'd184; b = 8'd163;  #10 
a = 8'd184; b = 8'd164;  #10 
a = 8'd184; b = 8'd165;  #10 
a = 8'd184; b = 8'd166;  #10 
a = 8'd184; b = 8'd167;  #10 
a = 8'd184; b = 8'd168;  #10 
a = 8'd184; b = 8'd169;  #10 
a = 8'd184; b = 8'd170;  #10 
a = 8'd184; b = 8'd171;  #10 
a = 8'd184; b = 8'd172;  #10 
a = 8'd184; b = 8'd173;  #10 
a = 8'd184; b = 8'd174;  #10 
a = 8'd184; b = 8'd175;  #10 
a = 8'd184; b = 8'd176;  #10 
a = 8'd184; b = 8'd177;  #10 
a = 8'd184; b = 8'd178;  #10 
a = 8'd184; b = 8'd179;  #10 
a = 8'd184; b = 8'd180;  #10 
a = 8'd184; b = 8'd181;  #10 
a = 8'd184; b = 8'd182;  #10 
a = 8'd184; b = 8'd183;  #10 
a = 8'd184; b = 8'd184;  #10 
a = 8'd184; b = 8'd185;  #10 
a = 8'd184; b = 8'd186;  #10 
a = 8'd184; b = 8'd187;  #10 
a = 8'd184; b = 8'd188;  #10 
a = 8'd184; b = 8'd189;  #10 
a = 8'd184; b = 8'd190;  #10 
a = 8'd184; b = 8'd191;  #10 
a = 8'd184; b = 8'd192;  #10 
a = 8'd184; b = 8'd193;  #10 
a = 8'd184; b = 8'd194;  #10 
a = 8'd184; b = 8'd195;  #10 
a = 8'd184; b = 8'd196;  #10 
a = 8'd184; b = 8'd197;  #10 
a = 8'd184; b = 8'd198;  #10 
a = 8'd184; b = 8'd199;  #10 
a = 8'd184; b = 8'd200;  #10 
a = 8'd184; b = 8'd201;  #10 
a = 8'd184; b = 8'd202;  #10 
a = 8'd184; b = 8'd203;  #10 
a = 8'd184; b = 8'd204;  #10 
a = 8'd184; b = 8'd205;  #10 
a = 8'd184; b = 8'd206;  #10 
a = 8'd184; b = 8'd207;  #10 
a = 8'd184; b = 8'd208;  #10 
a = 8'd184; b = 8'd209;  #10 
a = 8'd184; b = 8'd210;  #10 
a = 8'd184; b = 8'd211;  #10 
a = 8'd184; b = 8'd212;  #10 
a = 8'd184; b = 8'd213;  #10 
a = 8'd184; b = 8'd214;  #10 
a = 8'd184; b = 8'd215;  #10 
a = 8'd184; b = 8'd216;  #10 
a = 8'd184; b = 8'd217;  #10 
a = 8'd184; b = 8'd218;  #10 
a = 8'd184; b = 8'd219;  #10 
a = 8'd184; b = 8'd220;  #10 
a = 8'd184; b = 8'd221;  #10 
a = 8'd184; b = 8'd222;  #10 
a = 8'd184; b = 8'd223;  #10 
a = 8'd184; b = 8'd224;  #10 
a = 8'd184; b = 8'd225;  #10 
a = 8'd184; b = 8'd226;  #10 
a = 8'd184; b = 8'd227;  #10 
a = 8'd184; b = 8'd228;  #10 
a = 8'd184; b = 8'd229;  #10 
a = 8'd184; b = 8'd230;  #10 
a = 8'd184; b = 8'd231;  #10 
a = 8'd184; b = 8'd232;  #10 
a = 8'd184; b = 8'd233;  #10 
a = 8'd184; b = 8'd234;  #10 
a = 8'd184; b = 8'd235;  #10 
a = 8'd184; b = 8'd236;  #10 
a = 8'd184; b = 8'd237;  #10 
a = 8'd184; b = 8'd238;  #10 
a = 8'd184; b = 8'd239;  #10 
a = 8'd184; b = 8'd240;  #10 
a = 8'd184; b = 8'd241;  #10 
a = 8'd184; b = 8'd242;  #10 
a = 8'd184; b = 8'd243;  #10 
a = 8'd184; b = 8'd244;  #10 
a = 8'd184; b = 8'd245;  #10 
a = 8'd184; b = 8'd246;  #10 
a = 8'd184; b = 8'd247;  #10 
a = 8'd184; b = 8'd248;  #10 
a = 8'd184; b = 8'd249;  #10 
a = 8'd184; b = 8'd250;  #10 
a = 8'd184; b = 8'd251;  #10 
a = 8'd184; b = 8'd252;  #10 
a = 8'd184; b = 8'd253;  #10 
a = 8'd184; b = 8'd254;  #10 
a = 8'd184; b = 8'd255;  #10 
a = 8'd185; b = 8'd0;  #10 
a = 8'd185; b = 8'd1;  #10 
a = 8'd185; b = 8'd2;  #10 
a = 8'd185; b = 8'd3;  #10 
a = 8'd185; b = 8'd4;  #10 
a = 8'd185; b = 8'd5;  #10 
a = 8'd185; b = 8'd6;  #10 
a = 8'd185; b = 8'd7;  #10 
a = 8'd185; b = 8'd8;  #10 
a = 8'd185; b = 8'd9;  #10 
a = 8'd185; b = 8'd10;  #10 
a = 8'd185; b = 8'd11;  #10 
a = 8'd185; b = 8'd12;  #10 
a = 8'd185; b = 8'd13;  #10 
a = 8'd185; b = 8'd14;  #10 
a = 8'd185; b = 8'd15;  #10 
a = 8'd185; b = 8'd16;  #10 
a = 8'd185; b = 8'd17;  #10 
a = 8'd185; b = 8'd18;  #10 
a = 8'd185; b = 8'd19;  #10 
a = 8'd185; b = 8'd20;  #10 
a = 8'd185; b = 8'd21;  #10 
a = 8'd185; b = 8'd22;  #10 
a = 8'd185; b = 8'd23;  #10 
a = 8'd185; b = 8'd24;  #10 
a = 8'd185; b = 8'd25;  #10 
a = 8'd185; b = 8'd26;  #10 
a = 8'd185; b = 8'd27;  #10 
a = 8'd185; b = 8'd28;  #10 
a = 8'd185; b = 8'd29;  #10 
a = 8'd185; b = 8'd30;  #10 
a = 8'd185; b = 8'd31;  #10 
a = 8'd185; b = 8'd32;  #10 
a = 8'd185; b = 8'd33;  #10 
a = 8'd185; b = 8'd34;  #10 
a = 8'd185; b = 8'd35;  #10 
a = 8'd185; b = 8'd36;  #10 
a = 8'd185; b = 8'd37;  #10 
a = 8'd185; b = 8'd38;  #10 
a = 8'd185; b = 8'd39;  #10 
a = 8'd185; b = 8'd40;  #10 
a = 8'd185; b = 8'd41;  #10 
a = 8'd185; b = 8'd42;  #10 
a = 8'd185; b = 8'd43;  #10 
a = 8'd185; b = 8'd44;  #10 
a = 8'd185; b = 8'd45;  #10 
a = 8'd185; b = 8'd46;  #10 
a = 8'd185; b = 8'd47;  #10 
a = 8'd185; b = 8'd48;  #10 
a = 8'd185; b = 8'd49;  #10 
a = 8'd185; b = 8'd50;  #10 
a = 8'd185; b = 8'd51;  #10 
a = 8'd185; b = 8'd52;  #10 
a = 8'd185; b = 8'd53;  #10 
a = 8'd185; b = 8'd54;  #10 
a = 8'd185; b = 8'd55;  #10 
a = 8'd185; b = 8'd56;  #10 
a = 8'd185; b = 8'd57;  #10 
a = 8'd185; b = 8'd58;  #10 
a = 8'd185; b = 8'd59;  #10 
a = 8'd185; b = 8'd60;  #10 
a = 8'd185; b = 8'd61;  #10 
a = 8'd185; b = 8'd62;  #10 
a = 8'd185; b = 8'd63;  #10 
a = 8'd185; b = 8'd64;  #10 
a = 8'd185; b = 8'd65;  #10 
a = 8'd185; b = 8'd66;  #10 
a = 8'd185; b = 8'd67;  #10 
a = 8'd185; b = 8'd68;  #10 
a = 8'd185; b = 8'd69;  #10 
a = 8'd185; b = 8'd70;  #10 
a = 8'd185; b = 8'd71;  #10 
a = 8'd185; b = 8'd72;  #10 
a = 8'd185; b = 8'd73;  #10 
a = 8'd185; b = 8'd74;  #10 
a = 8'd185; b = 8'd75;  #10 
a = 8'd185; b = 8'd76;  #10 
a = 8'd185; b = 8'd77;  #10 
a = 8'd185; b = 8'd78;  #10 
a = 8'd185; b = 8'd79;  #10 
a = 8'd185; b = 8'd80;  #10 
a = 8'd185; b = 8'd81;  #10 
a = 8'd185; b = 8'd82;  #10 
a = 8'd185; b = 8'd83;  #10 
a = 8'd185; b = 8'd84;  #10 
a = 8'd185; b = 8'd85;  #10 
a = 8'd185; b = 8'd86;  #10 
a = 8'd185; b = 8'd87;  #10 
a = 8'd185; b = 8'd88;  #10 
a = 8'd185; b = 8'd89;  #10 
a = 8'd185; b = 8'd90;  #10 
a = 8'd185; b = 8'd91;  #10 
a = 8'd185; b = 8'd92;  #10 
a = 8'd185; b = 8'd93;  #10 
a = 8'd185; b = 8'd94;  #10 
a = 8'd185; b = 8'd95;  #10 
a = 8'd185; b = 8'd96;  #10 
a = 8'd185; b = 8'd97;  #10 
a = 8'd185; b = 8'd98;  #10 
a = 8'd185; b = 8'd99;  #10 
a = 8'd185; b = 8'd100;  #10 
a = 8'd185; b = 8'd101;  #10 
a = 8'd185; b = 8'd102;  #10 
a = 8'd185; b = 8'd103;  #10 
a = 8'd185; b = 8'd104;  #10 
a = 8'd185; b = 8'd105;  #10 
a = 8'd185; b = 8'd106;  #10 
a = 8'd185; b = 8'd107;  #10 
a = 8'd185; b = 8'd108;  #10 
a = 8'd185; b = 8'd109;  #10 
a = 8'd185; b = 8'd110;  #10 
a = 8'd185; b = 8'd111;  #10 
a = 8'd185; b = 8'd112;  #10 
a = 8'd185; b = 8'd113;  #10 
a = 8'd185; b = 8'd114;  #10 
a = 8'd185; b = 8'd115;  #10 
a = 8'd185; b = 8'd116;  #10 
a = 8'd185; b = 8'd117;  #10 
a = 8'd185; b = 8'd118;  #10 
a = 8'd185; b = 8'd119;  #10 
a = 8'd185; b = 8'd120;  #10 
a = 8'd185; b = 8'd121;  #10 
a = 8'd185; b = 8'd122;  #10 
a = 8'd185; b = 8'd123;  #10 
a = 8'd185; b = 8'd124;  #10 
a = 8'd185; b = 8'd125;  #10 
a = 8'd185; b = 8'd126;  #10 
a = 8'd185; b = 8'd127;  #10 
a = 8'd185; b = 8'd128;  #10 
a = 8'd185; b = 8'd129;  #10 
a = 8'd185; b = 8'd130;  #10 
a = 8'd185; b = 8'd131;  #10 
a = 8'd185; b = 8'd132;  #10 
a = 8'd185; b = 8'd133;  #10 
a = 8'd185; b = 8'd134;  #10 
a = 8'd185; b = 8'd135;  #10 
a = 8'd185; b = 8'd136;  #10 
a = 8'd185; b = 8'd137;  #10 
a = 8'd185; b = 8'd138;  #10 
a = 8'd185; b = 8'd139;  #10 
a = 8'd185; b = 8'd140;  #10 
a = 8'd185; b = 8'd141;  #10 
a = 8'd185; b = 8'd142;  #10 
a = 8'd185; b = 8'd143;  #10 
a = 8'd185; b = 8'd144;  #10 
a = 8'd185; b = 8'd145;  #10 
a = 8'd185; b = 8'd146;  #10 
a = 8'd185; b = 8'd147;  #10 
a = 8'd185; b = 8'd148;  #10 
a = 8'd185; b = 8'd149;  #10 
a = 8'd185; b = 8'd150;  #10 
a = 8'd185; b = 8'd151;  #10 
a = 8'd185; b = 8'd152;  #10 
a = 8'd185; b = 8'd153;  #10 
a = 8'd185; b = 8'd154;  #10 
a = 8'd185; b = 8'd155;  #10 
a = 8'd185; b = 8'd156;  #10 
a = 8'd185; b = 8'd157;  #10 
a = 8'd185; b = 8'd158;  #10 
a = 8'd185; b = 8'd159;  #10 
a = 8'd185; b = 8'd160;  #10 
a = 8'd185; b = 8'd161;  #10 
a = 8'd185; b = 8'd162;  #10 
a = 8'd185; b = 8'd163;  #10 
a = 8'd185; b = 8'd164;  #10 
a = 8'd185; b = 8'd165;  #10 
a = 8'd185; b = 8'd166;  #10 
a = 8'd185; b = 8'd167;  #10 
a = 8'd185; b = 8'd168;  #10 
a = 8'd185; b = 8'd169;  #10 
a = 8'd185; b = 8'd170;  #10 
a = 8'd185; b = 8'd171;  #10 
a = 8'd185; b = 8'd172;  #10 
a = 8'd185; b = 8'd173;  #10 
a = 8'd185; b = 8'd174;  #10 
a = 8'd185; b = 8'd175;  #10 
a = 8'd185; b = 8'd176;  #10 
a = 8'd185; b = 8'd177;  #10 
a = 8'd185; b = 8'd178;  #10 
a = 8'd185; b = 8'd179;  #10 
a = 8'd185; b = 8'd180;  #10 
a = 8'd185; b = 8'd181;  #10 
a = 8'd185; b = 8'd182;  #10 
a = 8'd185; b = 8'd183;  #10 
a = 8'd185; b = 8'd184;  #10 
a = 8'd185; b = 8'd185;  #10 
a = 8'd185; b = 8'd186;  #10 
a = 8'd185; b = 8'd187;  #10 
a = 8'd185; b = 8'd188;  #10 
a = 8'd185; b = 8'd189;  #10 
a = 8'd185; b = 8'd190;  #10 
a = 8'd185; b = 8'd191;  #10 
a = 8'd185; b = 8'd192;  #10 
a = 8'd185; b = 8'd193;  #10 
a = 8'd185; b = 8'd194;  #10 
a = 8'd185; b = 8'd195;  #10 
a = 8'd185; b = 8'd196;  #10 
a = 8'd185; b = 8'd197;  #10 
a = 8'd185; b = 8'd198;  #10 
a = 8'd185; b = 8'd199;  #10 
a = 8'd185; b = 8'd200;  #10 
a = 8'd185; b = 8'd201;  #10 
a = 8'd185; b = 8'd202;  #10 
a = 8'd185; b = 8'd203;  #10 
a = 8'd185; b = 8'd204;  #10 
a = 8'd185; b = 8'd205;  #10 
a = 8'd185; b = 8'd206;  #10 
a = 8'd185; b = 8'd207;  #10 
a = 8'd185; b = 8'd208;  #10 
a = 8'd185; b = 8'd209;  #10 
a = 8'd185; b = 8'd210;  #10 
a = 8'd185; b = 8'd211;  #10 
a = 8'd185; b = 8'd212;  #10 
a = 8'd185; b = 8'd213;  #10 
a = 8'd185; b = 8'd214;  #10 
a = 8'd185; b = 8'd215;  #10 
a = 8'd185; b = 8'd216;  #10 
a = 8'd185; b = 8'd217;  #10 
a = 8'd185; b = 8'd218;  #10 
a = 8'd185; b = 8'd219;  #10 
a = 8'd185; b = 8'd220;  #10 
a = 8'd185; b = 8'd221;  #10 
a = 8'd185; b = 8'd222;  #10 
a = 8'd185; b = 8'd223;  #10 
a = 8'd185; b = 8'd224;  #10 
a = 8'd185; b = 8'd225;  #10 
a = 8'd185; b = 8'd226;  #10 
a = 8'd185; b = 8'd227;  #10 
a = 8'd185; b = 8'd228;  #10 
a = 8'd185; b = 8'd229;  #10 
a = 8'd185; b = 8'd230;  #10 
a = 8'd185; b = 8'd231;  #10 
a = 8'd185; b = 8'd232;  #10 
a = 8'd185; b = 8'd233;  #10 
a = 8'd185; b = 8'd234;  #10 
a = 8'd185; b = 8'd235;  #10 
a = 8'd185; b = 8'd236;  #10 
a = 8'd185; b = 8'd237;  #10 
a = 8'd185; b = 8'd238;  #10 
a = 8'd185; b = 8'd239;  #10 
a = 8'd185; b = 8'd240;  #10 
a = 8'd185; b = 8'd241;  #10 
a = 8'd185; b = 8'd242;  #10 
a = 8'd185; b = 8'd243;  #10 
a = 8'd185; b = 8'd244;  #10 
a = 8'd185; b = 8'd245;  #10 
a = 8'd185; b = 8'd246;  #10 
a = 8'd185; b = 8'd247;  #10 
a = 8'd185; b = 8'd248;  #10 
a = 8'd185; b = 8'd249;  #10 
a = 8'd185; b = 8'd250;  #10 
a = 8'd185; b = 8'd251;  #10 
a = 8'd185; b = 8'd252;  #10 
a = 8'd185; b = 8'd253;  #10 
a = 8'd185; b = 8'd254;  #10 
a = 8'd185; b = 8'd255;  #10 
a = 8'd186; b = 8'd0;  #10 
a = 8'd186; b = 8'd1;  #10 
a = 8'd186; b = 8'd2;  #10 
a = 8'd186; b = 8'd3;  #10 
a = 8'd186; b = 8'd4;  #10 
a = 8'd186; b = 8'd5;  #10 
a = 8'd186; b = 8'd6;  #10 
a = 8'd186; b = 8'd7;  #10 
a = 8'd186; b = 8'd8;  #10 
a = 8'd186; b = 8'd9;  #10 
a = 8'd186; b = 8'd10;  #10 
a = 8'd186; b = 8'd11;  #10 
a = 8'd186; b = 8'd12;  #10 
a = 8'd186; b = 8'd13;  #10 
a = 8'd186; b = 8'd14;  #10 
a = 8'd186; b = 8'd15;  #10 
a = 8'd186; b = 8'd16;  #10 
a = 8'd186; b = 8'd17;  #10 
a = 8'd186; b = 8'd18;  #10 
a = 8'd186; b = 8'd19;  #10 
a = 8'd186; b = 8'd20;  #10 
a = 8'd186; b = 8'd21;  #10 
a = 8'd186; b = 8'd22;  #10 
a = 8'd186; b = 8'd23;  #10 
a = 8'd186; b = 8'd24;  #10 
a = 8'd186; b = 8'd25;  #10 
a = 8'd186; b = 8'd26;  #10 
a = 8'd186; b = 8'd27;  #10 
a = 8'd186; b = 8'd28;  #10 
a = 8'd186; b = 8'd29;  #10 
a = 8'd186; b = 8'd30;  #10 
a = 8'd186; b = 8'd31;  #10 
a = 8'd186; b = 8'd32;  #10 
a = 8'd186; b = 8'd33;  #10 
a = 8'd186; b = 8'd34;  #10 
a = 8'd186; b = 8'd35;  #10 
a = 8'd186; b = 8'd36;  #10 
a = 8'd186; b = 8'd37;  #10 
a = 8'd186; b = 8'd38;  #10 
a = 8'd186; b = 8'd39;  #10 
a = 8'd186; b = 8'd40;  #10 
a = 8'd186; b = 8'd41;  #10 
a = 8'd186; b = 8'd42;  #10 
a = 8'd186; b = 8'd43;  #10 
a = 8'd186; b = 8'd44;  #10 
a = 8'd186; b = 8'd45;  #10 
a = 8'd186; b = 8'd46;  #10 
a = 8'd186; b = 8'd47;  #10 
a = 8'd186; b = 8'd48;  #10 
a = 8'd186; b = 8'd49;  #10 
a = 8'd186; b = 8'd50;  #10 
a = 8'd186; b = 8'd51;  #10 
a = 8'd186; b = 8'd52;  #10 
a = 8'd186; b = 8'd53;  #10 
a = 8'd186; b = 8'd54;  #10 
a = 8'd186; b = 8'd55;  #10 
a = 8'd186; b = 8'd56;  #10 
a = 8'd186; b = 8'd57;  #10 
a = 8'd186; b = 8'd58;  #10 
a = 8'd186; b = 8'd59;  #10 
a = 8'd186; b = 8'd60;  #10 
a = 8'd186; b = 8'd61;  #10 
a = 8'd186; b = 8'd62;  #10 
a = 8'd186; b = 8'd63;  #10 
a = 8'd186; b = 8'd64;  #10 
a = 8'd186; b = 8'd65;  #10 
a = 8'd186; b = 8'd66;  #10 
a = 8'd186; b = 8'd67;  #10 
a = 8'd186; b = 8'd68;  #10 
a = 8'd186; b = 8'd69;  #10 
a = 8'd186; b = 8'd70;  #10 
a = 8'd186; b = 8'd71;  #10 
a = 8'd186; b = 8'd72;  #10 
a = 8'd186; b = 8'd73;  #10 
a = 8'd186; b = 8'd74;  #10 
a = 8'd186; b = 8'd75;  #10 
a = 8'd186; b = 8'd76;  #10 
a = 8'd186; b = 8'd77;  #10 
a = 8'd186; b = 8'd78;  #10 
a = 8'd186; b = 8'd79;  #10 
a = 8'd186; b = 8'd80;  #10 
a = 8'd186; b = 8'd81;  #10 
a = 8'd186; b = 8'd82;  #10 
a = 8'd186; b = 8'd83;  #10 
a = 8'd186; b = 8'd84;  #10 
a = 8'd186; b = 8'd85;  #10 
a = 8'd186; b = 8'd86;  #10 
a = 8'd186; b = 8'd87;  #10 
a = 8'd186; b = 8'd88;  #10 
a = 8'd186; b = 8'd89;  #10 
a = 8'd186; b = 8'd90;  #10 
a = 8'd186; b = 8'd91;  #10 
a = 8'd186; b = 8'd92;  #10 
a = 8'd186; b = 8'd93;  #10 
a = 8'd186; b = 8'd94;  #10 
a = 8'd186; b = 8'd95;  #10 
a = 8'd186; b = 8'd96;  #10 
a = 8'd186; b = 8'd97;  #10 
a = 8'd186; b = 8'd98;  #10 
a = 8'd186; b = 8'd99;  #10 
a = 8'd186; b = 8'd100;  #10 
a = 8'd186; b = 8'd101;  #10 
a = 8'd186; b = 8'd102;  #10 
a = 8'd186; b = 8'd103;  #10 
a = 8'd186; b = 8'd104;  #10 
a = 8'd186; b = 8'd105;  #10 
a = 8'd186; b = 8'd106;  #10 
a = 8'd186; b = 8'd107;  #10 
a = 8'd186; b = 8'd108;  #10 
a = 8'd186; b = 8'd109;  #10 
a = 8'd186; b = 8'd110;  #10 
a = 8'd186; b = 8'd111;  #10 
a = 8'd186; b = 8'd112;  #10 
a = 8'd186; b = 8'd113;  #10 
a = 8'd186; b = 8'd114;  #10 
a = 8'd186; b = 8'd115;  #10 
a = 8'd186; b = 8'd116;  #10 
a = 8'd186; b = 8'd117;  #10 
a = 8'd186; b = 8'd118;  #10 
a = 8'd186; b = 8'd119;  #10 
a = 8'd186; b = 8'd120;  #10 
a = 8'd186; b = 8'd121;  #10 
a = 8'd186; b = 8'd122;  #10 
a = 8'd186; b = 8'd123;  #10 
a = 8'd186; b = 8'd124;  #10 
a = 8'd186; b = 8'd125;  #10 
a = 8'd186; b = 8'd126;  #10 
a = 8'd186; b = 8'd127;  #10 
a = 8'd186; b = 8'd128;  #10 
a = 8'd186; b = 8'd129;  #10 
a = 8'd186; b = 8'd130;  #10 
a = 8'd186; b = 8'd131;  #10 
a = 8'd186; b = 8'd132;  #10 
a = 8'd186; b = 8'd133;  #10 
a = 8'd186; b = 8'd134;  #10 
a = 8'd186; b = 8'd135;  #10 
a = 8'd186; b = 8'd136;  #10 
a = 8'd186; b = 8'd137;  #10 
a = 8'd186; b = 8'd138;  #10 
a = 8'd186; b = 8'd139;  #10 
a = 8'd186; b = 8'd140;  #10 
a = 8'd186; b = 8'd141;  #10 
a = 8'd186; b = 8'd142;  #10 
a = 8'd186; b = 8'd143;  #10 
a = 8'd186; b = 8'd144;  #10 
a = 8'd186; b = 8'd145;  #10 
a = 8'd186; b = 8'd146;  #10 
a = 8'd186; b = 8'd147;  #10 
a = 8'd186; b = 8'd148;  #10 
a = 8'd186; b = 8'd149;  #10 
a = 8'd186; b = 8'd150;  #10 
a = 8'd186; b = 8'd151;  #10 
a = 8'd186; b = 8'd152;  #10 
a = 8'd186; b = 8'd153;  #10 
a = 8'd186; b = 8'd154;  #10 
a = 8'd186; b = 8'd155;  #10 
a = 8'd186; b = 8'd156;  #10 
a = 8'd186; b = 8'd157;  #10 
a = 8'd186; b = 8'd158;  #10 
a = 8'd186; b = 8'd159;  #10 
a = 8'd186; b = 8'd160;  #10 
a = 8'd186; b = 8'd161;  #10 
a = 8'd186; b = 8'd162;  #10 
a = 8'd186; b = 8'd163;  #10 
a = 8'd186; b = 8'd164;  #10 
a = 8'd186; b = 8'd165;  #10 
a = 8'd186; b = 8'd166;  #10 
a = 8'd186; b = 8'd167;  #10 
a = 8'd186; b = 8'd168;  #10 
a = 8'd186; b = 8'd169;  #10 
a = 8'd186; b = 8'd170;  #10 
a = 8'd186; b = 8'd171;  #10 
a = 8'd186; b = 8'd172;  #10 
a = 8'd186; b = 8'd173;  #10 
a = 8'd186; b = 8'd174;  #10 
a = 8'd186; b = 8'd175;  #10 
a = 8'd186; b = 8'd176;  #10 
a = 8'd186; b = 8'd177;  #10 
a = 8'd186; b = 8'd178;  #10 
a = 8'd186; b = 8'd179;  #10 
a = 8'd186; b = 8'd180;  #10 
a = 8'd186; b = 8'd181;  #10 
a = 8'd186; b = 8'd182;  #10 
a = 8'd186; b = 8'd183;  #10 
a = 8'd186; b = 8'd184;  #10 
a = 8'd186; b = 8'd185;  #10 
a = 8'd186; b = 8'd186;  #10 
a = 8'd186; b = 8'd187;  #10 
a = 8'd186; b = 8'd188;  #10 
a = 8'd186; b = 8'd189;  #10 
a = 8'd186; b = 8'd190;  #10 
a = 8'd186; b = 8'd191;  #10 
a = 8'd186; b = 8'd192;  #10 
a = 8'd186; b = 8'd193;  #10 
a = 8'd186; b = 8'd194;  #10 
a = 8'd186; b = 8'd195;  #10 
a = 8'd186; b = 8'd196;  #10 
a = 8'd186; b = 8'd197;  #10 
a = 8'd186; b = 8'd198;  #10 
a = 8'd186; b = 8'd199;  #10 
a = 8'd186; b = 8'd200;  #10 
a = 8'd186; b = 8'd201;  #10 
a = 8'd186; b = 8'd202;  #10 
a = 8'd186; b = 8'd203;  #10 
a = 8'd186; b = 8'd204;  #10 
a = 8'd186; b = 8'd205;  #10 
a = 8'd186; b = 8'd206;  #10 
a = 8'd186; b = 8'd207;  #10 
a = 8'd186; b = 8'd208;  #10 
a = 8'd186; b = 8'd209;  #10 
a = 8'd186; b = 8'd210;  #10 
a = 8'd186; b = 8'd211;  #10 
a = 8'd186; b = 8'd212;  #10 
a = 8'd186; b = 8'd213;  #10 
a = 8'd186; b = 8'd214;  #10 
a = 8'd186; b = 8'd215;  #10 
a = 8'd186; b = 8'd216;  #10 
a = 8'd186; b = 8'd217;  #10 
a = 8'd186; b = 8'd218;  #10 
a = 8'd186; b = 8'd219;  #10 
a = 8'd186; b = 8'd220;  #10 
a = 8'd186; b = 8'd221;  #10 
a = 8'd186; b = 8'd222;  #10 
a = 8'd186; b = 8'd223;  #10 
a = 8'd186; b = 8'd224;  #10 
a = 8'd186; b = 8'd225;  #10 
a = 8'd186; b = 8'd226;  #10 
a = 8'd186; b = 8'd227;  #10 
a = 8'd186; b = 8'd228;  #10 
a = 8'd186; b = 8'd229;  #10 
a = 8'd186; b = 8'd230;  #10 
a = 8'd186; b = 8'd231;  #10 
a = 8'd186; b = 8'd232;  #10 
a = 8'd186; b = 8'd233;  #10 
a = 8'd186; b = 8'd234;  #10 
a = 8'd186; b = 8'd235;  #10 
a = 8'd186; b = 8'd236;  #10 
a = 8'd186; b = 8'd237;  #10 
a = 8'd186; b = 8'd238;  #10 
a = 8'd186; b = 8'd239;  #10 
a = 8'd186; b = 8'd240;  #10 
a = 8'd186; b = 8'd241;  #10 
a = 8'd186; b = 8'd242;  #10 
a = 8'd186; b = 8'd243;  #10 
a = 8'd186; b = 8'd244;  #10 
a = 8'd186; b = 8'd245;  #10 
a = 8'd186; b = 8'd246;  #10 
a = 8'd186; b = 8'd247;  #10 
a = 8'd186; b = 8'd248;  #10 
a = 8'd186; b = 8'd249;  #10 
a = 8'd186; b = 8'd250;  #10 
a = 8'd186; b = 8'd251;  #10 
a = 8'd186; b = 8'd252;  #10 
a = 8'd186; b = 8'd253;  #10 
a = 8'd186; b = 8'd254;  #10 
a = 8'd186; b = 8'd255;  #10 
a = 8'd187; b = 8'd0;  #10 
a = 8'd187; b = 8'd1;  #10 
a = 8'd187; b = 8'd2;  #10 
a = 8'd187; b = 8'd3;  #10 
a = 8'd187; b = 8'd4;  #10 
a = 8'd187; b = 8'd5;  #10 
a = 8'd187; b = 8'd6;  #10 
a = 8'd187; b = 8'd7;  #10 
a = 8'd187; b = 8'd8;  #10 
a = 8'd187; b = 8'd9;  #10 
a = 8'd187; b = 8'd10;  #10 
a = 8'd187; b = 8'd11;  #10 
a = 8'd187; b = 8'd12;  #10 
a = 8'd187; b = 8'd13;  #10 
a = 8'd187; b = 8'd14;  #10 
a = 8'd187; b = 8'd15;  #10 
a = 8'd187; b = 8'd16;  #10 
a = 8'd187; b = 8'd17;  #10 
a = 8'd187; b = 8'd18;  #10 
a = 8'd187; b = 8'd19;  #10 
a = 8'd187; b = 8'd20;  #10 
a = 8'd187; b = 8'd21;  #10 
a = 8'd187; b = 8'd22;  #10 
a = 8'd187; b = 8'd23;  #10 
a = 8'd187; b = 8'd24;  #10 
a = 8'd187; b = 8'd25;  #10 
a = 8'd187; b = 8'd26;  #10 
a = 8'd187; b = 8'd27;  #10 
a = 8'd187; b = 8'd28;  #10 
a = 8'd187; b = 8'd29;  #10 
a = 8'd187; b = 8'd30;  #10 
a = 8'd187; b = 8'd31;  #10 
a = 8'd187; b = 8'd32;  #10 
a = 8'd187; b = 8'd33;  #10 
a = 8'd187; b = 8'd34;  #10 
a = 8'd187; b = 8'd35;  #10 
a = 8'd187; b = 8'd36;  #10 
a = 8'd187; b = 8'd37;  #10 
a = 8'd187; b = 8'd38;  #10 
a = 8'd187; b = 8'd39;  #10 
a = 8'd187; b = 8'd40;  #10 
a = 8'd187; b = 8'd41;  #10 
a = 8'd187; b = 8'd42;  #10 
a = 8'd187; b = 8'd43;  #10 
a = 8'd187; b = 8'd44;  #10 
a = 8'd187; b = 8'd45;  #10 
a = 8'd187; b = 8'd46;  #10 
a = 8'd187; b = 8'd47;  #10 
a = 8'd187; b = 8'd48;  #10 
a = 8'd187; b = 8'd49;  #10 
a = 8'd187; b = 8'd50;  #10 
a = 8'd187; b = 8'd51;  #10 
a = 8'd187; b = 8'd52;  #10 
a = 8'd187; b = 8'd53;  #10 
a = 8'd187; b = 8'd54;  #10 
a = 8'd187; b = 8'd55;  #10 
a = 8'd187; b = 8'd56;  #10 
a = 8'd187; b = 8'd57;  #10 
a = 8'd187; b = 8'd58;  #10 
a = 8'd187; b = 8'd59;  #10 
a = 8'd187; b = 8'd60;  #10 
a = 8'd187; b = 8'd61;  #10 
a = 8'd187; b = 8'd62;  #10 
a = 8'd187; b = 8'd63;  #10 
a = 8'd187; b = 8'd64;  #10 
a = 8'd187; b = 8'd65;  #10 
a = 8'd187; b = 8'd66;  #10 
a = 8'd187; b = 8'd67;  #10 
a = 8'd187; b = 8'd68;  #10 
a = 8'd187; b = 8'd69;  #10 
a = 8'd187; b = 8'd70;  #10 
a = 8'd187; b = 8'd71;  #10 
a = 8'd187; b = 8'd72;  #10 
a = 8'd187; b = 8'd73;  #10 
a = 8'd187; b = 8'd74;  #10 
a = 8'd187; b = 8'd75;  #10 
a = 8'd187; b = 8'd76;  #10 
a = 8'd187; b = 8'd77;  #10 
a = 8'd187; b = 8'd78;  #10 
a = 8'd187; b = 8'd79;  #10 
a = 8'd187; b = 8'd80;  #10 
a = 8'd187; b = 8'd81;  #10 
a = 8'd187; b = 8'd82;  #10 
a = 8'd187; b = 8'd83;  #10 
a = 8'd187; b = 8'd84;  #10 
a = 8'd187; b = 8'd85;  #10 
a = 8'd187; b = 8'd86;  #10 
a = 8'd187; b = 8'd87;  #10 
a = 8'd187; b = 8'd88;  #10 
a = 8'd187; b = 8'd89;  #10 
a = 8'd187; b = 8'd90;  #10 
a = 8'd187; b = 8'd91;  #10 
a = 8'd187; b = 8'd92;  #10 
a = 8'd187; b = 8'd93;  #10 
a = 8'd187; b = 8'd94;  #10 
a = 8'd187; b = 8'd95;  #10 
a = 8'd187; b = 8'd96;  #10 
a = 8'd187; b = 8'd97;  #10 
a = 8'd187; b = 8'd98;  #10 
a = 8'd187; b = 8'd99;  #10 
a = 8'd187; b = 8'd100;  #10 
a = 8'd187; b = 8'd101;  #10 
a = 8'd187; b = 8'd102;  #10 
a = 8'd187; b = 8'd103;  #10 
a = 8'd187; b = 8'd104;  #10 
a = 8'd187; b = 8'd105;  #10 
a = 8'd187; b = 8'd106;  #10 
a = 8'd187; b = 8'd107;  #10 
a = 8'd187; b = 8'd108;  #10 
a = 8'd187; b = 8'd109;  #10 
a = 8'd187; b = 8'd110;  #10 
a = 8'd187; b = 8'd111;  #10 
a = 8'd187; b = 8'd112;  #10 
a = 8'd187; b = 8'd113;  #10 
a = 8'd187; b = 8'd114;  #10 
a = 8'd187; b = 8'd115;  #10 
a = 8'd187; b = 8'd116;  #10 
a = 8'd187; b = 8'd117;  #10 
a = 8'd187; b = 8'd118;  #10 
a = 8'd187; b = 8'd119;  #10 
a = 8'd187; b = 8'd120;  #10 
a = 8'd187; b = 8'd121;  #10 
a = 8'd187; b = 8'd122;  #10 
a = 8'd187; b = 8'd123;  #10 
a = 8'd187; b = 8'd124;  #10 
a = 8'd187; b = 8'd125;  #10 
a = 8'd187; b = 8'd126;  #10 
a = 8'd187; b = 8'd127;  #10 
a = 8'd187; b = 8'd128;  #10 
a = 8'd187; b = 8'd129;  #10 
a = 8'd187; b = 8'd130;  #10 
a = 8'd187; b = 8'd131;  #10 
a = 8'd187; b = 8'd132;  #10 
a = 8'd187; b = 8'd133;  #10 
a = 8'd187; b = 8'd134;  #10 
a = 8'd187; b = 8'd135;  #10 
a = 8'd187; b = 8'd136;  #10 
a = 8'd187; b = 8'd137;  #10 
a = 8'd187; b = 8'd138;  #10 
a = 8'd187; b = 8'd139;  #10 
a = 8'd187; b = 8'd140;  #10 
a = 8'd187; b = 8'd141;  #10 
a = 8'd187; b = 8'd142;  #10 
a = 8'd187; b = 8'd143;  #10 
a = 8'd187; b = 8'd144;  #10 
a = 8'd187; b = 8'd145;  #10 
a = 8'd187; b = 8'd146;  #10 
a = 8'd187; b = 8'd147;  #10 
a = 8'd187; b = 8'd148;  #10 
a = 8'd187; b = 8'd149;  #10 
a = 8'd187; b = 8'd150;  #10 
a = 8'd187; b = 8'd151;  #10 
a = 8'd187; b = 8'd152;  #10 
a = 8'd187; b = 8'd153;  #10 
a = 8'd187; b = 8'd154;  #10 
a = 8'd187; b = 8'd155;  #10 
a = 8'd187; b = 8'd156;  #10 
a = 8'd187; b = 8'd157;  #10 
a = 8'd187; b = 8'd158;  #10 
a = 8'd187; b = 8'd159;  #10 
a = 8'd187; b = 8'd160;  #10 
a = 8'd187; b = 8'd161;  #10 
a = 8'd187; b = 8'd162;  #10 
a = 8'd187; b = 8'd163;  #10 
a = 8'd187; b = 8'd164;  #10 
a = 8'd187; b = 8'd165;  #10 
a = 8'd187; b = 8'd166;  #10 
a = 8'd187; b = 8'd167;  #10 
a = 8'd187; b = 8'd168;  #10 
a = 8'd187; b = 8'd169;  #10 
a = 8'd187; b = 8'd170;  #10 
a = 8'd187; b = 8'd171;  #10 
a = 8'd187; b = 8'd172;  #10 
a = 8'd187; b = 8'd173;  #10 
a = 8'd187; b = 8'd174;  #10 
a = 8'd187; b = 8'd175;  #10 
a = 8'd187; b = 8'd176;  #10 
a = 8'd187; b = 8'd177;  #10 
a = 8'd187; b = 8'd178;  #10 
a = 8'd187; b = 8'd179;  #10 
a = 8'd187; b = 8'd180;  #10 
a = 8'd187; b = 8'd181;  #10 
a = 8'd187; b = 8'd182;  #10 
a = 8'd187; b = 8'd183;  #10 
a = 8'd187; b = 8'd184;  #10 
a = 8'd187; b = 8'd185;  #10 
a = 8'd187; b = 8'd186;  #10 
a = 8'd187; b = 8'd187;  #10 
a = 8'd187; b = 8'd188;  #10 
a = 8'd187; b = 8'd189;  #10 
a = 8'd187; b = 8'd190;  #10 
a = 8'd187; b = 8'd191;  #10 
a = 8'd187; b = 8'd192;  #10 
a = 8'd187; b = 8'd193;  #10 
a = 8'd187; b = 8'd194;  #10 
a = 8'd187; b = 8'd195;  #10 
a = 8'd187; b = 8'd196;  #10 
a = 8'd187; b = 8'd197;  #10 
a = 8'd187; b = 8'd198;  #10 
a = 8'd187; b = 8'd199;  #10 
a = 8'd187; b = 8'd200;  #10 
a = 8'd187; b = 8'd201;  #10 
a = 8'd187; b = 8'd202;  #10 
a = 8'd187; b = 8'd203;  #10 
a = 8'd187; b = 8'd204;  #10 
a = 8'd187; b = 8'd205;  #10 
a = 8'd187; b = 8'd206;  #10 
a = 8'd187; b = 8'd207;  #10 
a = 8'd187; b = 8'd208;  #10 
a = 8'd187; b = 8'd209;  #10 
a = 8'd187; b = 8'd210;  #10 
a = 8'd187; b = 8'd211;  #10 
a = 8'd187; b = 8'd212;  #10 
a = 8'd187; b = 8'd213;  #10 
a = 8'd187; b = 8'd214;  #10 
a = 8'd187; b = 8'd215;  #10 
a = 8'd187; b = 8'd216;  #10 
a = 8'd187; b = 8'd217;  #10 
a = 8'd187; b = 8'd218;  #10 
a = 8'd187; b = 8'd219;  #10 
a = 8'd187; b = 8'd220;  #10 
a = 8'd187; b = 8'd221;  #10 
a = 8'd187; b = 8'd222;  #10 
a = 8'd187; b = 8'd223;  #10 
a = 8'd187; b = 8'd224;  #10 
a = 8'd187; b = 8'd225;  #10 
a = 8'd187; b = 8'd226;  #10 
a = 8'd187; b = 8'd227;  #10 
a = 8'd187; b = 8'd228;  #10 
a = 8'd187; b = 8'd229;  #10 
a = 8'd187; b = 8'd230;  #10 
a = 8'd187; b = 8'd231;  #10 
a = 8'd187; b = 8'd232;  #10 
a = 8'd187; b = 8'd233;  #10 
a = 8'd187; b = 8'd234;  #10 
a = 8'd187; b = 8'd235;  #10 
a = 8'd187; b = 8'd236;  #10 
a = 8'd187; b = 8'd237;  #10 
a = 8'd187; b = 8'd238;  #10 
a = 8'd187; b = 8'd239;  #10 
a = 8'd187; b = 8'd240;  #10 
a = 8'd187; b = 8'd241;  #10 
a = 8'd187; b = 8'd242;  #10 
a = 8'd187; b = 8'd243;  #10 
a = 8'd187; b = 8'd244;  #10 
a = 8'd187; b = 8'd245;  #10 
a = 8'd187; b = 8'd246;  #10 
a = 8'd187; b = 8'd247;  #10 
a = 8'd187; b = 8'd248;  #10 
a = 8'd187; b = 8'd249;  #10 
a = 8'd187; b = 8'd250;  #10 
a = 8'd187; b = 8'd251;  #10 
a = 8'd187; b = 8'd252;  #10 
a = 8'd187; b = 8'd253;  #10 
a = 8'd187; b = 8'd254;  #10 
a = 8'd187; b = 8'd255;  #10 
a = 8'd188; b = 8'd0;  #10 
a = 8'd188; b = 8'd1;  #10 
a = 8'd188; b = 8'd2;  #10 
a = 8'd188; b = 8'd3;  #10 
a = 8'd188; b = 8'd4;  #10 
a = 8'd188; b = 8'd5;  #10 
a = 8'd188; b = 8'd6;  #10 
a = 8'd188; b = 8'd7;  #10 
a = 8'd188; b = 8'd8;  #10 
a = 8'd188; b = 8'd9;  #10 
a = 8'd188; b = 8'd10;  #10 
a = 8'd188; b = 8'd11;  #10 
a = 8'd188; b = 8'd12;  #10 
a = 8'd188; b = 8'd13;  #10 
a = 8'd188; b = 8'd14;  #10 
a = 8'd188; b = 8'd15;  #10 
a = 8'd188; b = 8'd16;  #10 
a = 8'd188; b = 8'd17;  #10 
a = 8'd188; b = 8'd18;  #10 
a = 8'd188; b = 8'd19;  #10 
a = 8'd188; b = 8'd20;  #10 
a = 8'd188; b = 8'd21;  #10 
a = 8'd188; b = 8'd22;  #10 
a = 8'd188; b = 8'd23;  #10 
a = 8'd188; b = 8'd24;  #10 
a = 8'd188; b = 8'd25;  #10 
a = 8'd188; b = 8'd26;  #10 
a = 8'd188; b = 8'd27;  #10 
a = 8'd188; b = 8'd28;  #10 
a = 8'd188; b = 8'd29;  #10 
a = 8'd188; b = 8'd30;  #10 
a = 8'd188; b = 8'd31;  #10 
a = 8'd188; b = 8'd32;  #10 
a = 8'd188; b = 8'd33;  #10 
a = 8'd188; b = 8'd34;  #10 
a = 8'd188; b = 8'd35;  #10 
a = 8'd188; b = 8'd36;  #10 
a = 8'd188; b = 8'd37;  #10 
a = 8'd188; b = 8'd38;  #10 
a = 8'd188; b = 8'd39;  #10 
a = 8'd188; b = 8'd40;  #10 
a = 8'd188; b = 8'd41;  #10 
a = 8'd188; b = 8'd42;  #10 
a = 8'd188; b = 8'd43;  #10 
a = 8'd188; b = 8'd44;  #10 
a = 8'd188; b = 8'd45;  #10 
a = 8'd188; b = 8'd46;  #10 
a = 8'd188; b = 8'd47;  #10 
a = 8'd188; b = 8'd48;  #10 
a = 8'd188; b = 8'd49;  #10 
a = 8'd188; b = 8'd50;  #10 
a = 8'd188; b = 8'd51;  #10 
a = 8'd188; b = 8'd52;  #10 
a = 8'd188; b = 8'd53;  #10 
a = 8'd188; b = 8'd54;  #10 
a = 8'd188; b = 8'd55;  #10 
a = 8'd188; b = 8'd56;  #10 
a = 8'd188; b = 8'd57;  #10 
a = 8'd188; b = 8'd58;  #10 
a = 8'd188; b = 8'd59;  #10 
a = 8'd188; b = 8'd60;  #10 
a = 8'd188; b = 8'd61;  #10 
a = 8'd188; b = 8'd62;  #10 
a = 8'd188; b = 8'd63;  #10 
a = 8'd188; b = 8'd64;  #10 
a = 8'd188; b = 8'd65;  #10 
a = 8'd188; b = 8'd66;  #10 
a = 8'd188; b = 8'd67;  #10 
a = 8'd188; b = 8'd68;  #10 
a = 8'd188; b = 8'd69;  #10 
a = 8'd188; b = 8'd70;  #10 
a = 8'd188; b = 8'd71;  #10 
a = 8'd188; b = 8'd72;  #10 
a = 8'd188; b = 8'd73;  #10 
a = 8'd188; b = 8'd74;  #10 
a = 8'd188; b = 8'd75;  #10 
a = 8'd188; b = 8'd76;  #10 
a = 8'd188; b = 8'd77;  #10 
a = 8'd188; b = 8'd78;  #10 
a = 8'd188; b = 8'd79;  #10 
a = 8'd188; b = 8'd80;  #10 
a = 8'd188; b = 8'd81;  #10 
a = 8'd188; b = 8'd82;  #10 
a = 8'd188; b = 8'd83;  #10 
a = 8'd188; b = 8'd84;  #10 
a = 8'd188; b = 8'd85;  #10 
a = 8'd188; b = 8'd86;  #10 
a = 8'd188; b = 8'd87;  #10 
a = 8'd188; b = 8'd88;  #10 
a = 8'd188; b = 8'd89;  #10 
a = 8'd188; b = 8'd90;  #10 
a = 8'd188; b = 8'd91;  #10 
a = 8'd188; b = 8'd92;  #10 
a = 8'd188; b = 8'd93;  #10 
a = 8'd188; b = 8'd94;  #10 
a = 8'd188; b = 8'd95;  #10 
a = 8'd188; b = 8'd96;  #10 
a = 8'd188; b = 8'd97;  #10 
a = 8'd188; b = 8'd98;  #10 
a = 8'd188; b = 8'd99;  #10 
a = 8'd188; b = 8'd100;  #10 
a = 8'd188; b = 8'd101;  #10 
a = 8'd188; b = 8'd102;  #10 
a = 8'd188; b = 8'd103;  #10 
a = 8'd188; b = 8'd104;  #10 
a = 8'd188; b = 8'd105;  #10 
a = 8'd188; b = 8'd106;  #10 
a = 8'd188; b = 8'd107;  #10 
a = 8'd188; b = 8'd108;  #10 
a = 8'd188; b = 8'd109;  #10 
a = 8'd188; b = 8'd110;  #10 
a = 8'd188; b = 8'd111;  #10 
a = 8'd188; b = 8'd112;  #10 
a = 8'd188; b = 8'd113;  #10 
a = 8'd188; b = 8'd114;  #10 
a = 8'd188; b = 8'd115;  #10 
a = 8'd188; b = 8'd116;  #10 
a = 8'd188; b = 8'd117;  #10 
a = 8'd188; b = 8'd118;  #10 
a = 8'd188; b = 8'd119;  #10 
a = 8'd188; b = 8'd120;  #10 
a = 8'd188; b = 8'd121;  #10 
a = 8'd188; b = 8'd122;  #10 
a = 8'd188; b = 8'd123;  #10 
a = 8'd188; b = 8'd124;  #10 
a = 8'd188; b = 8'd125;  #10 
a = 8'd188; b = 8'd126;  #10 
a = 8'd188; b = 8'd127;  #10 
a = 8'd188; b = 8'd128;  #10 
a = 8'd188; b = 8'd129;  #10 
a = 8'd188; b = 8'd130;  #10 
a = 8'd188; b = 8'd131;  #10 
a = 8'd188; b = 8'd132;  #10 
a = 8'd188; b = 8'd133;  #10 
a = 8'd188; b = 8'd134;  #10 
a = 8'd188; b = 8'd135;  #10 
a = 8'd188; b = 8'd136;  #10 
a = 8'd188; b = 8'd137;  #10 
a = 8'd188; b = 8'd138;  #10 
a = 8'd188; b = 8'd139;  #10 
a = 8'd188; b = 8'd140;  #10 
a = 8'd188; b = 8'd141;  #10 
a = 8'd188; b = 8'd142;  #10 
a = 8'd188; b = 8'd143;  #10 
a = 8'd188; b = 8'd144;  #10 
a = 8'd188; b = 8'd145;  #10 
a = 8'd188; b = 8'd146;  #10 
a = 8'd188; b = 8'd147;  #10 
a = 8'd188; b = 8'd148;  #10 
a = 8'd188; b = 8'd149;  #10 
a = 8'd188; b = 8'd150;  #10 
a = 8'd188; b = 8'd151;  #10 
a = 8'd188; b = 8'd152;  #10 
a = 8'd188; b = 8'd153;  #10 
a = 8'd188; b = 8'd154;  #10 
a = 8'd188; b = 8'd155;  #10 
a = 8'd188; b = 8'd156;  #10 
a = 8'd188; b = 8'd157;  #10 
a = 8'd188; b = 8'd158;  #10 
a = 8'd188; b = 8'd159;  #10 
a = 8'd188; b = 8'd160;  #10 
a = 8'd188; b = 8'd161;  #10 
a = 8'd188; b = 8'd162;  #10 
a = 8'd188; b = 8'd163;  #10 
a = 8'd188; b = 8'd164;  #10 
a = 8'd188; b = 8'd165;  #10 
a = 8'd188; b = 8'd166;  #10 
a = 8'd188; b = 8'd167;  #10 
a = 8'd188; b = 8'd168;  #10 
a = 8'd188; b = 8'd169;  #10 
a = 8'd188; b = 8'd170;  #10 
a = 8'd188; b = 8'd171;  #10 
a = 8'd188; b = 8'd172;  #10 
a = 8'd188; b = 8'd173;  #10 
a = 8'd188; b = 8'd174;  #10 
a = 8'd188; b = 8'd175;  #10 
a = 8'd188; b = 8'd176;  #10 
a = 8'd188; b = 8'd177;  #10 
a = 8'd188; b = 8'd178;  #10 
a = 8'd188; b = 8'd179;  #10 
a = 8'd188; b = 8'd180;  #10 
a = 8'd188; b = 8'd181;  #10 
a = 8'd188; b = 8'd182;  #10 
a = 8'd188; b = 8'd183;  #10 
a = 8'd188; b = 8'd184;  #10 
a = 8'd188; b = 8'd185;  #10 
a = 8'd188; b = 8'd186;  #10 
a = 8'd188; b = 8'd187;  #10 
a = 8'd188; b = 8'd188;  #10 
a = 8'd188; b = 8'd189;  #10 
a = 8'd188; b = 8'd190;  #10 
a = 8'd188; b = 8'd191;  #10 
a = 8'd188; b = 8'd192;  #10 
a = 8'd188; b = 8'd193;  #10 
a = 8'd188; b = 8'd194;  #10 
a = 8'd188; b = 8'd195;  #10 
a = 8'd188; b = 8'd196;  #10 
a = 8'd188; b = 8'd197;  #10 
a = 8'd188; b = 8'd198;  #10 
a = 8'd188; b = 8'd199;  #10 
a = 8'd188; b = 8'd200;  #10 
a = 8'd188; b = 8'd201;  #10 
a = 8'd188; b = 8'd202;  #10 
a = 8'd188; b = 8'd203;  #10 
a = 8'd188; b = 8'd204;  #10 
a = 8'd188; b = 8'd205;  #10 
a = 8'd188; b = 8'd206;  #10 
a = 8'd188; b = 8'd207;  #10 
a = 8'd188; b = 8'd208;  #10 
a = 8'd188; b = 8'd209;  #10 
a = 8'd188; b = 8'd210;  #10 
a = 8'd188; b = 8'd211;  #10 
a = 8'd188; b = 8'd212;  #10 
a = 8'd188; b = 8'd213;  #10 
a = 8'd188; b = 8'd214;  #10 
a = 8'd188; b = 8'd215;  #10 
a = 8'd188; b = 8'd216;  #10 
a = 8'd188; b = 8'd217;  #10 
a = 8'd188; b = 8'd218;  #10 
a = 8'd188; b = 8'd219;  #10 
a = 8'd188; b = 8'd220;  #10 
a = 8'd188; b = 8'd221;  #10 
a = 8'd188; b = 8'd222;  #10 
a = 8'd188; b = 8'd223;  #10 
a = 8'd188; b = 8'd224;  #10 
a = 8'd188; b = 8'd225;  #10 
a = 8'd188; b = 8'd226;  #10 
a = 8'd188; b = 8'd227;  #10 
a = 8'd188; b = 8'd228;  #10 
a = 8'd188; b = 8'd229;  #10 
a = 8'd188; b = 8'd230;  #10 
a = 8'd188; b = 8'd231;  #10 
a = 8'd188; b = 8'd232;  #10 
a = 8'd188; b = 8'd233;  #10 
a = 8'd188; b = 8'd234;  #10 
a = 8'd188; b = 8'd235;  #10 
a = 8'd188; b = 8'd236;  #10 
a = 8'd188; b = 8'd237;  #10 
a = 8'd188; b = 8'd238;  #10 
a = 8'd188; b = 8'd239;  #10 
a = 8'd188; b = 8'd240;  #10 
a = 8'd188; b = 8'd241;  #10 
a = 8'd188; b = 8'd242;  #10 
a = 8'd188; b = 8'd243;  #10 
a = 8'd188; b = 8'd244;  #10 
a = 8'd188; b = 8'd245;  #10 
a = 8'd188; b = 8'd246;  #10 
a = 8'd188; b = 8'd247;  #10 
a = 8'd188; b = 8'd248;  #10 
a = 8'd188; b = 8'd249;  #10 
a = 8'd188; b = 8'd250;  #10 
a = 8'd188; b = 8'd251;  #10 
a = 8'd188; b = 8'd252;  #10 
a = 8'd188; b = 8'd253;  #10 
a = 8'd188; b = 8'd254;  #10 
a = 8'd188; b = 8'd255;  #10 
a = 8'd189; b = 8'd0;  #10 
a = 8'd189; b = 8'd1;  #10 
a = 8'd189; b = 8'd2;  #10 
a = 8'd189; b = 8'd3;  #10 
a = 8'd189; b = 8'd4;  #10 
a = 8'd189; b = 8'd5;  #10 
a = 8'd189; b = 8'd6;  #10 
a = 8'd189; b = 8'd7;  #10 
a = 8'd189; b = 8'd8;  #10 
a = 8'd189; b = 8'd9;  #10 
a = 8'd189; b = 8'd10;  #10 
a = 8'd189; b = 8'd11;  #10 
a = 8'd189; b = 8'd12;  #10 
a = 8'd189; b = 8'd13;  #10 
a = 8'd189; b = 8'd14;  #10 
a = 8'd189; b = 8'd15;  #10 
a = 8'd189; b = 8'd16;  #10 
a = 8'd189; b = 8'd17;  #10 
a = 8'd189; b = 8'd18;  #10 
a = 8'd189; b = 8'd19;  #10 
a = 8'd189; b = 8'd20;  #10 
a = 8'd189; b = 8'd21;  #10 
a = 8'd189; b = 8'd22;  #10 
a = 8'd189; b = 8'd23;  #10 
a = 8'd189; b = 8'd24;  #10 
a = 8'd189; b = 8'd25;  #10 
a = 8'd189; b = 8'd26;  #10 
a = 8'd189; b = 8'd27;  #10 
a = 8'd189; b = 8'd28;  #10 
a = 8'd189; b = 8'd29;  #10 
a = 8'd189; b = 8'd30;  #10 
a = 8'd189; b = 8'd31;  #10 
a = 8'd189; b = 8'd32;  #10 
a = 8'd189; b = 8'd33;  #10 
a = 8'd189; b = 8'd34;  #10 
a = 8'd189; b = 8'd35;  #10 
a = 8'd189; b = 8'd36;  #10 
a = 8'd189; b = 8'd37;  #10 
a = 8'd189; b = 8'd38;  #10 
a = 8'd189; b = 8'd39;  #10 
a = 8'd189; b = 8'd40;  #10 
a = 8'd189; b = 8'd41;  #10 
a = 8'd189; b = 8'd42;  #10 
a = 8'd189; b = 8'd43;  #10 
a = 8'd189; b = 8'd44;  #10 
a = 8'd189; b = 8'd45;  #10 
a = 8'd189; b = 8'd46;  #10 
a = 8'd189; b = 8'd47;  #10 
a = 8'd189; b = 8'd48;  #10 
a = 8'd189; b = 8'd49;  #10 
a = 8'd189; b = 8'd50;  #10 
a = 8'd189; b = 8'd51;  #10 
a = 8'd189; b = 8'd52;  #10 
a = 8'd189; b = 8'd53;  #10 
a = 8'd189; b = 8'd54;  #10 
a = 8'd189; b = 8'd55;  #10 
a = 8'd189; b = 8'd56;  #10 
a = 8'd189; b = 8'd57;  #10 
a = 8'd189; b = 8'd58;  #10 
a = 8'd189; b = 8'd59;  #10 
a = 8'd189; b = 8'd60;  #10 
a = 8'd189; b = 8'd61;  #10 
a = 8'd189; b = 8'd62;  #10 
a = 8'd189; b = 8'd63;  #10 
a = 8'd189; b = 8'd64;  #10 
a = 8'd189; b = 8'd65;  #10 
a = 8'd189; b = 8'd66;  #10 
a = 8'd189; b = 8'd67;  #10 
a = 8'd189; b = 8'd68;  #10 
a = 8'd189; b = 8'd69;  #10 
a = 8'd189; b = 8'd70;  #10 
a = 8'd189; b = 8'd71;  #10 
a = 8'd189; b = 8'd72;  #10 
a = 8'd189; b = 8'd73;  #10 
a = 8'd189; b = 8'd74;  #10 
a = 8'd189; b = 8'd75;  #10 
a = 8'd189; b = 8'd76;  #10 
a = 8'd189; b = 8'd77;  #10 
a = 8'd189; b = 8'd78;  #10 
a = 8'd189; b = 8'd79;  #10 
a = 8'd189; b = 8'd80;  #10 
a = 8'd189; b = 8'd81;  #10 
a = 8'd189; b = 8'd82;  #10 
a = 8'd189; b = 8'd83;  #10 
a = 8'd189; b = 8'd84;  #10 
a = 8'd189; b = 8'd85;  #10 
a = 8'd189; b = 8'd86;  #10 
a = 8'd189; b = 8'd87;  #10 
a = 8'd189; b = 8'd88;  #10 
a = 8'd189; b = 8'd89;  #10 
a = 8'd189; b = 8'd90;  #10 
a = 8'd189; b = 8'd91;  #10 
a = 8'd189; b = 8'd92;  #10 
a = 8'd189; b = 8'd93;  #10 
a = 8'd189; b = 8'd94;  #10 
a = 8'd189; b = 8'd95;  #10 
a = 8'd189; b = 8'd96;  #10 
a = 8'd189; b = 8'd97;  #10 
a = 8'd189; b = 8'd98;  #10 
a = 8'd189; b = 8'd99;  #10 
a = 8'd189; b = 8'd100;  #10 
a = 8'd189; b = 8'd101;  #10 
a = 8'd189; b = 8'd102;  #10 
a = 8'd189; b = 8'd103;  #10 
a = 8'd189; b = 8'd104;  #10 
a = 8'd189; b = 8'd105;  #10 
a = 8'd189; b = 8'd106;  #10 
a = 8'd189; b = 8'd107;  #10 
a = 8'd189; b = 8'd108;  #10 
a = 8'd189; b = 8'd109;  #10 
a = 8'd189; b = 8'd110;  #10 
a = 8'd189; b = 8'd111;  #10 
a = 8'd189; b = 8'd112;  #10 
a = 8'd189; b = 8'd113;  #10 
a = 8'd189; b = 8'd114;  #10 
a = 8'd189; b = 8'd115;  #10 
a = 8'd189; b = 8'd116;  #10 
a = 8'd189; b = 8'd117;  #10 
a = 8'd189; b = 8'd118;  #10 
a = 8'd189; b = 8'd119;  #10 
a = 8'd189; b = 8'd120;  #10 
a = 8'd189; b = 8'd121;  #10 
a = 8'd189; b = 8'd122;  #10 
a = 8'd189; b = 8'd123;  #10 
a = 8'd189; b = 8'd124;  #10 
a = 8'd189; b = 8'd125;  #10 
a = 8'd189; b = 8'd126;  #10 
a = 8'd189; b = 8'd127;  #10 
a = 8'd189; b = 8'd128;  #10 
a = 8'd189; b = 8'd129;  #10 
a = 8'd189; b = 8'd130;  #10 
a = 8'd189; b = 8'd131;  #10 
a = 8'd189; b = 8'd132;  #10 
a = 8'd189; b = 8'd133;  #10 
a = 8'd189; b = 8'd134;  #10 
a = 8'd189; b = 8'd135;  #10 
a = 8'd189; b = 8'd136;  #10 
a = 8'd189; b = 8'd137;  #10 
a = 8'd189; b = 8'd138;  #10 
a = 8'd189; b = 8'd139;  #10 
a = 8'd189; b = 8'd140;  #10 
a = 8'd189; b = 8'd141;  #10 
a = 8'd189; b = 8'd142;  #10 
a = 8'd189; b = 8'd143;  #10 
a = 8'd189; b = 8'd144;  #10 
a = 8'd189; b = 8'd145;  #10 
a = 8'd189; b = 8'd146;  #10 
a = 8'd189; b = 8'd147;  #10 
a = 8'd189; b = 8'd148;  #10 
a = 8'd189; b = 8'd149;  #10 
a = 8'd189; b = 8'd150;  #10 
a = 8'd189; b = 8'd151;  #10 
a = 8'd189; b = 8'd152;  #10 
a = 8'd189; b = 8'd153;  #10 
a = 8'd189; b = 8'd154;  #10 
a = 8'd189; b = 8'd155;  #10 
a = 8'd189; b = 8'd156;  #10 
a = 8'd189; b = 8'd157;  #10 
a = 8'd189; b = 8'd158;  #10 
a = 8'd189; b = 8'd159;  #10 
a = 8'd189; b = 8'd160;  #10 
a = 8'd189; b = 8'd161;  #10 
a = 8'd189; b = 8'd162;  #10 
a = 8'd189; b = 8'd163;  #10 
a = 8'd189; b = 8'd164;  #10 
a = 8'd189; b = 8'd165;  #10 
a = 8'd189; b = 8'd166;  #10 
a = 8'd189; b = 8'd167;  #10 
a = 8'd189; b = 8'd168;  #10 
a = 8'd189; b = 8'd169;  #10 
a = 8'd189; b = 8'd170;  #10 
a = 8'd189; b = 8'd171;  #10 
a = 8'd189; b = 8'd172;  #10 
a = 8'd189; b = 8'd173;  #10 
a = 8'd189; b = 8'd174;  #10 
a = 8'd189; b = 8'd175;  #10 
a = 8'd189; b = 8'd176;  #10 
a = 8'd189; b = 8'd177;  #10 
a = 8'd189; b = 8'd178;  #10 
a = 8'd189; b = 8'd179;  #10 
a = 8'd189; b = 8'd180;  #10 
a = 8'd189; b = 8'd181;  #10 
a = 8'd189; b = 8'd182;  #10 
a = 8'd189; b = 8'd183;  #10 
a = 8'd189; b = 8'd184;  #10 
a = 8'd189; b = 8'd185;  #10 
a = 8'd189; b = 8'd186;  #10 
a = 8'd189; b = 8'd187;  #10 
a = 8'd189; b = 8'd188;  #10 
a = 8'd189; b = 8'd189;  #10 
a = 8'd189; b = 8'd190;  #10 
a = 8'd189; b = 8'd191;  #10 
a = 8'd189; b = 8'd192;  #10 
a = 8'd189; b = 8'd193;  #10 
a = 8'd189; b = 8'd194;  #10 
a = 8'd189; b = 8'd195;  #10 
a = 8'd189; b = 8'd196;  #10 
a = 8'd189; b = 8'd197;  #10 
a = 8'd189; b = 8'd198;  #10 
a = 8'd189; b = 8'd199;  #10 
a = 8'd189; b = 8'd200;  #10 
a = 8'd189; b = 8'd201;  #10 
a = 8'd189; b = 8'd202;  #10 
a = 8'd189; b = 8'd203;  #10 
a = 8'd189; b = 8'd204;  #10 
a = 8'd189; b = 8'd205;  #10 
a = 8'd189; b = 8'd206;  #10 
a = 8'd189; b = 8'd207;  #10 
a = 8'd189; b = 8'd208;  #10 
a = 8'd189; b = 8'd209;  #10 
a = 8'd189; b = 8'd210;  #10 
a = 8'd189; b = 8'd211;  #10 
a = 8'd189; b = 8'd212;  #10 
a = 8'd189; b = 8'd213;  #10 
a = 8'd189; b = 8'd214;  #10 
a = 8'd189; b = 8'd215;  #10 
a = 8'd189; b = 8'd216;  #10 
a = 8'd189; b = 8'd217;  #10 
a = 8'd189; b = 8'd218;  #10 
a = 8'd189; b = 8'd219;  #10 
a = 8'd189; b = 8'd220;  #10 
a = 8'd189; b = 8'd221;  #10 
a = 8'd189; b = 8'd222;  #10 
a = 8'd189; b = 8'd223;  #10 
a = 8'd189; b = 8'd224;  #10 
a = 8'd189; b = 8'd225;  #10 
a = 8'd189; b = 8'd226;  #10 
a = 8'd189; b = 8'd227;  #10 
a = 8'd189; b = 8'd228;  #10 
a = 8'd189; b = 8'd229;  #10 
a = 8'd189; b = 8'd230;  #10 
a = 8'd189; b = 8'd231;  #10 
a = 8'd189; b = 8'd232;  #10 
a = 8'd189; b = 8'd233;  #10 
a = 8'd189; b = 8'd234;  #10 
a = 8'd189; b = 8'd235;  #10 
a = 8'd189; b = 8'd236;  #10 
a = 8'd189; b = 8'd237;  #10 
a = 8'd189; b = 8'd238;  #10 
a = 8'd189; b = 8'd239;  #10 
a = 8'd189; b = 8'd240;  #10 
a = 8'd189; b = 8'd241;  #10 
a = 8'd189; b = 8'd242;  #10 
a = 8'd189; b = 8'd243;  #10 
a = 8'd189; b = 8'd244;  #10 
a = 8'd189; b = 8'd245;  #10 
a = 8'd189; b = 8'd246;  #10 
a = 8'd189; b = 8'd247;  #10 
a = 8'd189; b = 8'd248;  #10 
a = 8'd189; b = 8'd249;  #10 
a = 8'd189; b = 8'd250;  #10 
a = 8'd189; b = 8'd251;  #10 
a = 8'd189; b = 8'd252;  #10 
a = 8'd189; b = 8'd253;  #10 
a = 8'd189; b = 8'd254;  #10 
a = 8'd189; b = 8'd255;  #10 
a = 8'd190; b = 8'd0;  #10 
a = 8'd190; b = 8'd1;  #10 
a = 8'd190; b = 8'd2;  #10 
a = 8'd190; b = 8'd3;  #10 
a = 8'd190; b = 8'd4;  #10 
a = 8'd190; b = 8'd5;  #10 
a = 8'd190; b = 8'd6;  #10 
a = 8'd190; b = 8'd7;  #10 
a = 8'd190; b = 8'd8;  #10 
a = 8'd190; b = 8'd9;  #10 
a = 8'd190; b = 8'd10;  #10 
a = 8'd190; b = 8'd11;  #10 
a = 8'd190; b = 8'd12;  #10 
a = 8'd190; b = 8'd13;  #10 
a = 8'd190; b = 8'd14;  #10 
a = 8'd190; b = 8'd15;  #10 
a = 8'd190; b = 8'd16;  #10 
a = 8'd190; b = 8'd17;  #10 
a = 8'd190; b = 8'd18;  #10 
a = 8'd190; b = 8'd19;  #10 
a = 8'd190; b = 8'd20;  #10 
a = 8'd190; b = 8'd21;  #10 
a = 8'd190; b = 8'd22;  #10 
a = 8'd190; b = 8'd23;  #10 
a = 8'd190; b = 8'd24;  #10 
a = 8'd190; b = 8'd25;  #10 
a = 8'd190; b = 8'd26;  #10 
a = 8'd190; b = 8'd27;  #10 
a = 8'd190; b = 8'd28;  #10 
a = 8'd190; b = 8'd29;  #10 
a = 8'd190; b = 8'd30;  #10 
a = 8'd190; b = 8'd31;  #10 
a = 8'd190; b = 8'd32;  #10 
a = 8'd190; b = 8'd33;  #10 
a = 8'd190; b = 8'd34;  #10 
a = 8'd190; b = 8'd35;  #10 
a = 8'd190; b = 8'd36;  #10 
a = 8'd190; b = 8'd37;  #10 
a = 8'd190; b = 8'd38;  #10 
a = 8'd190; b = 8'd39;  #10 
a = 8'd190; b = 8'd40;  #10 
a = 8'd190; b = 8'd41;  #10 
a = 8'd190; b = 8'd42;  #10 
a = 8'd190; b = 8'd43;  #10 
a = 8'd190; b = 8'd44;  #10 
a = 8'd190; b = 8'd45;  #10 
a = 8'd190; b = 8'd46;  #10 
a = 8'd190; b = 8'd47;  #10 
a = 8'd190; b = 8'd48;  #10 
a = 8'd190; b = 8'd49;  #10 
a = 8'd190; b = 8'd50;  #10 
a = 8'd190; b = 8'd51;  #10 
a = 8'd190; b = 8'd52;  #10 
a = 8'd190; b = 8'd53;  #10 
a = 8'd190; b = 8'd54;  #10 
a = 8'd190; b = 8'd55;  #10 
a = 8'd190; b = 8'd56;  #10 
a = 8'd190; b = 8'd57;  #10 
a = 8'd190; b = 8'd58;  #10 
a = 8'd190; b = 8'd59;  #10 
a = 8'd190; b = 8'd60;  #10 
a = 8'd190; b = 8'd61;  #10 
a = 8'd190; b = 8'd62;  #10 
a = 8'd190; b = 8'd63;  #10 
a = 8'd190; b = 8'd64;  #10 
a = 8'd190; b = 8'd65;  #10 
a = 8'd190; b = 8'd66;  #10 
a = 8'd190; b = 8'd67;  #10 
a = 8'd190; b = 8'd68;  #10 
a = 8'd190; b = 8'd69;  #10 
a = 8'd190; b = 8'd70;  #10 
a = 8'd190; b = 8'd71;  #10 
a = 8'd190; b = 8'd72;  #10 
a = 8'd190; b = 8'd73;  #10 
a = 8'd190; b = 8'd74;  #10 
a = 8'd190; b = 8'd75;  #10 
a = 8'd190; b = 8'd76;  #10 
a = 8'd190; b = 8'd77;  #10 
a = 8'd190; b = 8'd78;  #10 
a = 8'd190; b = 8'd79;  #10 
a = 8'd190; b = 8'd80;  #10 
a = 8'd190; b = 8'd81;  #10 
a = 8'd190; b = 8'd82;  #10 
a = 8'd190; b = 8'd83;  #10 
a = 8'd190; b = 8'd84;  #10 
a = 8'd190; b = 8'd85;  #10 
a = 8'd190; b = 8'd86;  #10 
a = 8'd190; b = 8'd87;  #10 
a = 8'd190; b = 8'd88;  #10 
a = 8'd190; b = 8'd89;  #10 
a = 8'd190; b = 8'd90;  #10 
a = 8'd190; b = 8'd91;  #10 
a = 8'd190; b = 8'd92;  #10 
a = 8'd190; b = 8'd93;  #10 
a = 8'd190; b = 8'd94;  #10 
a = 8'd190; b = 8'd95;  #10 
a = 8'd190; b = 8'd96;  #10 
a = 8'd190; b = 8'd97;  #10 
a = 8'd190; b = 8'd98;  #10 
a = 8'd190; b = 8'd99;  #10 
a = 8'd190; b = 8'd100;  #10 
a = 8'd190; b = 8'd101;  #10 
a = 8'd190; b = 8'd102;  #10 
a = 8'd190; b = 8'd103;  #10 
a = 8'd190; b = 8'd104;  #10 
a = 8'd190; b = 8'd105;  #10 
a = 8'd190; b = 8'd106;  #10 
a = 8'd190; b = 8'd107;  #10 
a = 8'd190; b = 8'd108;  #10 
a = 8'd190; b = 8'd109;  #10 
a = 8'd190; b = 8'd110;  #10 
a = 8'd190; b = 8'd111;  #10 
a = 8'd190; b = 8'd112;  #10 
a = 8'd190; b = 8'd113;  #10 
a = 8'd190; b = 8'd114;  #10 
a = 8'd190; b = 8'd115;  #10 
a = 8'd190; b = 8'd116;  #10 
a = 8'd190; b = 8'd117;  #10 
a = 8'd190; b = 8'd118;  #10 
a = 8'd190; b = 8'd119;  #10 
a = 8'd190; b = 8'd120;  #10 
a = 8'd190; b = 8'd121;  #10 
a = 8'd190; b = 8'd122;  #10 
a = 8'd190; b = 8'd123;  #10 
a = 8'd190; b = 8'd124;  #10 
a = 8'd190; b = 8'd125;  #10 
a = 8'd190; b = 8'd126;  #10 
a = 8'd190; b = 8'd127;  #10 
a = 8'd190; b = 8'd128;  #10 
a = 8'd190; b = 8'd129;  #10 
a = 8'd190; b = 8'd130;  #10 
a = 8'd190; b = 8'd131;  #10 
a = 8'd190; b = 8'd132;  #10 
a = 8'd190; b = 8'd133;  #10 
a = 8'd190; b = 8'd134;  #10 
a = 8'd190; b = 8'd135;  #10 
a = 8'd190; b = 8'd136;  #10 
a = 8'd190; b = 8'd137;  #10 
a = 8'd190; b = 8'd138;  #10 
a = 8'd190; b = 8'd139;  #10 
a = 8'd190; b = 8'd140;  #10 
a = 8'd190; b = 8'd141;  #10 
a = 8'd190; b = 8'd142;  #10 
a = 8'd190; b = 8'd143;  #10 
a = 8'd190; b = 8'd144;  #10 
a = 8'd190; b = 8'd145;  #10 
a = 8'd190; b = 8'd146;  #10 
a = 8'd190; b = 8'd147;  #10 
a = 8'd190; b = 8'd148;  #10 
a = 8'd190; b = 8'd149;  #10 
a = 8'd190; b = 8'd150;  #10 
a = 8'd190; b = 8'd151;  #10 
a = 8'd190; b = 8'd152;  #10 
a = 8'd190; b = 8'd153;  #10 
a = 8'd190; b = 8'd154;  #10 
a = 8'd190; b = 8'd155;  #10 
a = 8'd190; b = 8'd156;  #10 
a = 8'd190; b = 8'd157;  #10 
a = 8'd190; b = 8'd158;  #10 
a = 8'd190; b = 8'd159;  #10 
a = 8'd190; b = 8'd160;  #10 
a = 8'd190; b = 8'd161;  #10 
a = 8'd190; b = 8'd162;  #10 
a = 8'd190; b = 8'd163;  #10 
a = 8'd190; b = 8'd164;  #10 
a = 8'd190; b = 8'd165;  #10 
a = 8'd190; b = 8'd166;  #10 
a = 8'd190; b = 8'd167;  #10 
a = 8'd190; b = 8'd168;  #10 
a = 8'd190; b = 8'd169;  #10 
a = 8'd190; b = 8'd170;  #10 
a = 8'd190; b = 8'd171;  #10 
a = 8'd190; b = 8'd172;  #10 
a = 8'd190; b = 8'd173;  #10 
a = 8'd190; b = 8'd174;  #10 
a = 8'd190; b = 8'd175;  #10 
a = 8'd190; b = 8'd176;  #10 
a = 8'd190; b = 8'd177;  #10 
a = 8'd190; b = 8'd178;  #10 
a = 8'd190; b = 8'd179;  #10 
a = 8'd190; b = 8'd180;  #10 
a = 8'd190; b = 8'd181;  #10 
a = 8'd190; b = 8'd182;  #10 
a = 8'd190; b = 8'd183;  #10 
a = 8'd190; b = 8'd184;  #10 
a = 8'd190; b = 8'd185;  #10 
a = 8'd190; b = 8'd186;  #10 
a = 8'd190; b = 8'd187;  #10 
a = 8'd190; b = 8'd188;  #10 
a = 8'd190; b = 8'd189;  #10 
a = 8'd190; b = 8'd190;  #10 
a = 8'd190; b = 8'd191;  #10 
a = 8'd190; b = 8'd192;  #10 
a = 8'd190; b = 8'd193;  #10 
a = 8'd190; b = 8'd194;  #10 
a = 8'd190; b = 8'd195;  #10 
a = 8'd190; b = 8'd196;  #10 
a = 8'd190; b = 8'd197;  #10 
a = 8'd190; b = 8'd198;  #10 
a = 8'd190; b = 8'd199;  #10 
a = 8'd190; b = 8'd200;  #10 
a = 8'd190; b = 8'd201;  #10 
a = 8'd190; b = 8'd202;  #10 
a = 8'd190; b = 8'd203;  #10 
a = 8'd190; b = 8'd204;  #10 
a = 8'd190; b = 8'd205;  #10 
a = 8'd190; b = 8'd206;  #10 
a = 8'd190; b = 8'd207;  #10 
a = 8'd190; b = 8'd208;  #10 
a = 8'd190; b = 8'd209;  #10 
a = 8'd190; b = 8'd210;  #10 
a = 8'd190; b = 8'd211;  #10 
a = 8'd190; b = 8'd212;  #10 
a = 8'd190; b = 8'd213;  #10 
a = 8'd190; b = 8'd214;  #10 
a = 8'd190; b = 8'd215;  #10 
a = 8'd190; b = 8'd216;  #10 
a = 8'd190; b = 8'd217;  #10 
a = 8'd190; b = 8'd218;  #10 
a = 8'd190; b = 8'd219;  #10 
a = 8'd190; b = 8'd220;  #10 
a = 8'd190; b = 8'd221;  #10 
a = 8'd190; b = 8'd222;  #10 
a = 8'd190; b = 8'd223;  #10 
a = 8'd190; b = 8'd224;  #10 
a = 8'd190; b = 8'd225;  #10 
a = 8'd190; b = 8'd226;  #10 
a = 8'd190; b = 8'd227;  #10 
a = 8'd190; b = 8'd228;  #10 
a = 8'd190; b = 8'd229;  #10 
a = 8'd190; b = 8'd230;  #10 
a = 8'd190; b = 8'd231;  #10 
a = 8'd190; b = 8'd232;  #10 
a = 8'd190; b = 8'd233;  #10 
a = 8'd190; b = 8'd234;  #10 
a = 8'd190; b = 8'd235;  #10 
a = 8'd190; b = 8'd236;  #10 
a = 8'd190; b = 8'd237;  #10 
a = 8'd190; b = 8'd238;  #10 
a = 8'd190; b = 8'd239;  #10 
a = 8'd190; b = 8'd240;  #10 
a = 8'd190; b = 8'd241;  #10 
a = 8'd190; b = 8'd242;  #10 
a = 8'd190; b = 8'd243;  #10 
a = 8'd190; b = 8'd244;  #10 
a = 8'd190; b = 8'd245;  #10 
a = 8'd190; b = 8'd246;  #10 
a = 8'd190; b = 8'd247;  #10 
a = 8'd190; b = 8'd248;  #10 
a = 8'd190; b = 8'd249;  #10 
a = 8'd190; b = 8'd250;  #10 
a = 8'd190; b = 8'd251;  #10 
a = 8'd190; b = 8'd252;  #10 
a = 8'd190; b = 8'd253;  #10 
a = 8'd190; b = 8'd254;  #10 
a = 8'd190; b = 8'd255;  #10 
a = 8'd191; b = 8'd0;  #10 
a = 8'd191; b = 8'd1;  #10 
a = 8'd191; b = 8'd2;  #10 
a = 8'd191; b = 8'd3;  #10 
a = 8'd191; b = 8'd4;  #10 
a = 8'd191; b = 8'd5;  #10 
a = 8'd191; b = 8'd6;  #10 
a = 8'd191; b = 8'd7;  #10 
a = 8'd191; b = 8'd8;  #10 
a = 8'd191; b = 8'd9;  #10 
a = 8'd191; b = 8'd10;  #10 
a = 8'd191; b = 8'd11;  #10 
a = 8'd191; b = 8'd12;  #10 
a = 8'd191; b = 8'd13;  #10 
a = 8'd191; b = 8'd14;  #10 
a = 8'd191; b = 8'd15;  #10 
a = 8'd191; b = 8'd16;  #10 
a = 8'd191; b = 8'd17;  #10 
a = 8'd191; b = 8'd18;  #10 
a = 8'd191; b = 8'd19;  #10 
a = 8'd191; b = 8'd20;  #10 
a = 8'd191; b = 8'd21;  #10 
a = 8'd191; b = 8'd22;  #10 
a = 8'd191; b = 8'd23;  #10 
a = 8'd191; b = 8'd24;  #10 
a = 8'd191; b = 8'd25;  #10 
a = 8'd191; b = 8'd26;  #10 
a = 8'd191; b = 8'd27;  #10 
a = 8'd191; b = 8'd28;  #10 
a = 8'd191; b = 8'd29;  #10 
a = 8'd191; b = 8'd30;  #10 
a = 8'd191; b = 8'd31;  #10 
a = 8'd191; b = 8'd32;  #10 
a = 8'd191; b = 8'd33;  #10 
a = 8'd191; b = 8'd34;  #10 
a = 8'd191; b = 8'd35;  #10 
a = 8'd191; b = 8'd36;  #10 
a = 8'd191; b = 8'd37;  #10 
a = 8'd191; b = 8'd38;  #10 
a = 8'd191; b = 8'd39;  #10 
a = 8'd191; b = 8'd40;  #10 
a = 8'd191; b = 8'd41;  #10 
a = 8'd191; b = 8'd42;  #10 
a = 8'd191; b = 8'd43;  #10 
a = 8'd191; b = 8'd44;  #10 
a = 8'd191; b = 8'd45;  #10 
a = 8'd191; b = 8'd46;  #10 
a = 8'd191; b = 8'd47;  #10 
a = 8'd191; b = 8'd48;  #10 
a = 8'd191; b = 8'd49;  #10 
a = 8'd191; b = 8'd50;  #10 
a = 8'd191; b = 8'd51;  #10 
a = 8'd191; b = 8'd52;  #10 
a = 8'd191; b = 8'd53;  #10 
a = 8'd191; b = 8'd54;  #10 
a = 8'd191; b = 8'd55;  #10 
a = 8'd191; b = 8'd56;  #10 
a = 8'd191; b = 8'd57;  #10 
a = 8'd191; b = 8'd58;  #10 
a = 8'd191; b = 8'd59;  #10 
a = 8'd191; b = 8'd60;  #10 
a = 8'd191; b = 8'd61;  #10 
a = 8'd191; b = 8'd62;  #10 
a = 8'd191; b = 8'd63;  #10 
a = 8'd191; b = 8'd64;  #10 
a = 8'd191; b = 8'd65;  #10 
a = 8'd191; b = 8'd66;  #10 
a = 8'd191; b = 8'd67;  #10 
a = 8'd191; b = 8'd68;  #10 
a = 8'd191; b = 8'd69;  #10 
a = 8'd191; b = 8'd70;  #10 
a = 8'd191; b = 8'd71;  #10 
a = 8'd191; b = 8'd72;  #10 
a = 8'd191; b = 8'd73;  #10 
a = 8'd191; b = 8'd74;  #10 
a = 8'd191; b = 8'd75;  #10 
a = 8'd191; b = 8'd76;  #10 
a = 8'd191; b = 8'd77;  #10 
a = 8'd191; b = 8'd78;  #10 
a = 8'd191; b = 8'd79;  #10 
a = 8'd191; b = 8'd80;  #10 
a = 8'd191; b = 8'd81;  #10 
a = 8'd191; b = 8'd82;  #10 
a = 8'd191; b = 8'd83;  #10 
a = 8'd191; b = 8'd84;  #10 
a = 8'd191; b = 8'd85;  #10 
a = 8'd191; b = 8'd86;  #10 
a = 8'd191; b = 8'd87;  #10 
a = 8'd191; b = 8'd88;  #10 
a = 8'd191; b = 8'd89;  #10 
a = 8'd191; b = 8'd90;  #10 
a = 8'd191; b = 8'd91;  #10 
a = 8'd191; b = 8'd92;  #10 
a = 8'd191; b = 8'd93;  #10 
a = 8'd191; b = 8'd94;  #10 
a = 8'd191; b = 8'd95;  #10 
a = 8'd191; b = 8'd96;  #10 
a = 8'd191; b = 8'd97;  #10 
a = 8'd191; b = 8'd98;  #10 
a = 8'd191; b = 8'd99;  #10 
a = 8'd191; b = 8'd100;  #10 
a = 8'd191; b = 8'd101;  #10 
a = 8'd191; b = 8'd102;  #10 
a = 8'd191; b = 8'd103;  #10 
a = 8'd191; b = 8'd104;  #10 
a = 8'd191; b = 8'd105;  #10 
a = 8'd191; b = 8'd106;  #10 
a = 8'd191; b = 8'd107;  #10 
a = 8'd191; b = 8'd108;  #10 
a = 8'd191; b = 8'd109;  #10 
a = 8'd191; b = 8'd110;  #10 
a = 8'd191; b = 8'd111;  #10 
a = 8'd191; b = 8'd112;  #10 
a = 8'd191; b = 8'd113;  #10 
a = 8'd191; b = 8'd114;  #10 
a = 8'd191; b = 8'd115;  #10 
a = 8'd191; b = 8'd116;  #10 
a = 8'd191; b = 8'd117;  #10 
a = 8'd191; b = 8'd118;  #10 
a = 8'd191; b = 8'd119;  #10 
a = 8'd191; b = 8'd120;  #10 
a = 8'd191; b = 8'd121;  #10 
a = 8'd191; b = 8'd122;  #10 
a = 8'd191; b = 8'd123;  #10 
a = 8'd191; b = 8'd124;  #10 
a = 8'd191; b = 8'd125;  #10 
a = 8'd191; b = 8'd126;  #10 
a = 8'd191; b = 8'd127;  #10 
a = 8'd191; b = 8'd128;  #10 
a = 8'd191; b = 8'd129;  #10 
a = 8'd191; b = 8'd130;  #10 
a = 8'd191; b = 8'd131;  #10 
a = 8'd191; b = 8'd132;  #10 
a = 8'd191; b = 8'd133;  #10 
a = 8'd191; b = 8'd134;  #10 
a = 8'd191; b = 8'd135;  #10 
a = 8'd191; b = 8'd136;  #10 
a = 8'd191; b = 8'd137;  #10 
a = 8'd191; b = 8'd138;  #10 
a = 8'd191; b = 8'd139;  #10 
a = 8'd191; b = 8'd140;  #10 
a = 8'd191; b = 8'd141;  #10 
a = 8'd191; b = 8'd142;  #10 
a = 8'd191; b = 8'd143;  #10 
a = 8'd191; b = 8'd144;  #10 
a = 8'd191; b = 8'd145;  #10 
a = 8'd191; b = 8'd146;  #10 
a = 8'd191; b = 8'd147;  #10 
a = 8'd191; b = 8'd148;  #10 
a = 8'd191; b = 8'd149;  #10 
a = 8'd191; b = 8'd150;  #10 
a = 8'd191; b = 8'd151;  #10 
a = 8'd191; b = 8'd152;  #10 
a = 8'd191; b = 8'd153;  #10 
a = 8'd191; b = 8'd154;  #10 
a = 8'd191; b = 8'd155;  #10 
a = 8'd191; b = 8'd156;  #10 
a = 8'd191; b = 8'd157;  #10 
a = 8'd191; b = 8'd158;  #10 
a = 8'd191; b = 8'd159;  #10 
a = 8'd191; b = 8'd160;  #10 
a = 8'd191; b = 8'd161;  #10 
a = 8'd191; b = 8'd162;  #10 
a = 8'd191; b = 8'd163;  #10 
a = 8'd191; b = 8'd164;  #10 
a = 8'd191; b = 8'd165;  #10 
a = 8'd191; b = 8'd166;  #10 
a = 8'd191; b = 8'd167;  #10 
a = 8'd191; b = 8'd168;  #10 
a = 8'd191; b = 8'd169;  #10 
a = 8'd191; b = 8'd170;  #10 
a = 8'd191; b = 8'd171;  #10 
a = 8'd191; b = 8'd172;  #10 
a = 8'd191; b = 8'd173;  #10 
a = 8'd191; b = 8'd174;  #10 
a = 8'd191; b = 8'd175;  #10 
a = 8'd191; b = 8'd176;  #10 
a = 8'd191; b = 8'd177;  #10 
a = 8'd191; b = 8'd178;  #10 
a = 8'd191; b = 8'd179;  #10 
a = 8'd191; b = 8'd180;  #10 
a = 8'd191; b = 8'd181;  #10 
a = 8'd191; b = 8'd182;  #10 
a = 8'd191; b = 8'd183;  #10 
a = 8'd191; b = 8'd184;  #10 
a = 8'd191; b = 8'd185;  #10 
a = 8'd191; b = 8'd186;  #10 
a = 8'd191; b = 8'd187;  #10 
a = 8'd191; b = 8'd188;  #10 
a = 8'd191; b = 8'd189;  #10 
a = 8'd191; b = 8'd190;  #10 
a = 8'd191; b = 8'd191;  #10 
a = 8'd191; b = 8'd192;  #10 
a = 8'd191; b = 8'd193;  #10 
a = 8'd191; b = 8'd194;  #10 
a = 8'd191; b = 8'd195;  #10 
a = 8'd191; b = 8'd196;  #10 
a = 8'd191; b = 8'd197;  #10 
a = 8'd191; b = 8'd198;  #10 
a = 8'd191; b = 8'd199;  #10 
a = 8'd191; b = 8'd200;  #10 
a = 8'd191; b = 8'd201;  #10 
a = 8'd191; b = 8'd202;  #10 
a = 8'd191; b = 8'd203;  #10 
a = 8'd191; b = 8'd204;  #10 
a = 8'd191; b = 8'd205;  #10 
a = 8'd191; b = 8'd206;  #10 
a = 8'd191; b = 8'd207;  #10 
a = 8'd191; b = 8'd208;  #10 
a = 8'd191; b = 8'd209;  #10 
a = 8'd191; b = 8'd210;  #10 
a = 8'd191; b = 8'd211;  #10 
a = 8'd191; b = 8'd212;  #10 
a = 8'd191; b = 8'd213;  #10 
a = 8'd191; b = 8'd214;  #10 
a = 8'd191; b = 8'd215;  #10 
a = 8'd191; b = 8'd216;  #10 
a = 8'd191; b = 8'd217;  #10 
a = 8'd191; b = 8'd218;  #10 
a = 8'd191; b = 8'd219;  #10 
a = 8'd191; b = 8'd220;  #10 
a = 8'd191; b = 8'd221;  #10 
a = 8'd191; b = 8'd222;  #10 
a = 8'd191; b = 8'd223;  #10 
a = 8'd191; b = 8'd224;  #10 
a = 8'd191; b = 8'd225;  #10 
a = 8'd191; b = 8'd226;  #10 
a = 8'd191; b = 8'd227;  #10 
a = 8'd191; b = 8'd228;  #10 
a = 8'd191; b = 8'd229;  #10 
a = 8'd191; b = 8'd230;  #10 
a = 8'd191; b = 8'd231;  #10 
a = 8'd191; b = 8'd232;  #10 
a = 8'd191; b = 8'd233;  #10 
a = 8'd191; b = 8'd234;  #10 
a = 8'd191; b = 8'd235;  #10 
a = 8'd191; b = 8'd236;  #10 
a = 8'd191; b = 8'd237;  #10 
a = 8'd191; b = 8'd238;  #10 
a = 8'd191; b = 8'd239;  #10 
a = 8'd191; b = 8'd240;  #10 
a = 8'd191; b = 8'd241;  #10 
a = 8'd191; b = 8'd242;  #10 
a = 8'd191; b = 8'd243;  #10 
a = 8'd191; b = 8'd244;  #10 
a = 8'd191; b = 8'd245;  #10 
a = 8'd191; b = 8'd246;  #10 
a = 8'd191; b = 8'd247;  #10 
a = 8'd191; b = 8'd248;  #10 
a = 8'd191; b = 8'd249;  #10 
a = 8'd191; b = 8'd250;  #10 
a = 8'd191; b = 8'd251;  #10 
a = 8'd191; b = 8'd252;  #10 
a = 8'd191; b = 8'd253;  #10 
a = 8'd191; b = 8'd254;  #10 
a = 8'd191; b = 8'd255;  #10 
a = 8'd192; b = 8'd0;  #10 
a = 8'd192; b = 8'd1;  #10 
a = 8'd192; b = 8'd2;  #10 
a = 8'd192; b = 8'd3;  #10 
a = 8'd192; b = 8'd4;  #10 
a = 8'd192; b = 8'd5;  #10 
a = 8'd192; b = 8'd6;  #10 
a = 8'd192; b = 8'd7;  #10 
a = 8'd192; b = 8'd8;  #10 
a = 8'd192; b = 8'd9;  #10 
a = 8'd192; b = 8'd10;  #10 
a = 8'd192; b = 8'd11;  #10 
a = 8'd192; b = 8'd12;  #10 
a = 8'd192; b = 8'd13;  #10 
a = 8'd192; b = 8'd14;  #10 
a = 8'd192; b = 8'd15;  #10 
a = 8'd192; b = 8'd16;  #10 
a = 8'd192; b = 8'd17;  #10 
a = 8'd192; b = 8'd18;  #10 
a = 8'd192; b = 8'd19;  #10 
a = 8'd192; b = 8'd20;  #10 
a = 8'd192; b = 8'd21;  #10 
a = 8'd192; b = 8'd22;  #10 
a = 8'd192; b = 8'd23;  #10 
a = 8'd192; b = 8'd24;  #10 
a = 8'd192; b = 8'd25;  #10 
a = 8'd192; b = 8'd26;  #10 
a = 8'd192; b = 8'd27;  #10 
a = 8'd192; b = 8'd28;  #10 
a = 8'd192; b = 8'd29;  #10 
a = 8'd192; b = 8'd30;  #10 
a = 8'd192; b = 8'd31;  #10 
a = 8'd192; b = 8'd32;  #10 
a = 8'd192; b = 8'd33;  #10 
a = 8'd192; b = 8'd34;  #10 
a = 8'd192; b = 8'd35;  #10 
a = 8'd192; b = 8'd36;  #10 
a = 8'd192; b = 8'd37;  #10 
a = 8'd192; b = 8'd38;  #10 
a = 8'd192; b = 8'd39;  #10 
a = 8'd192; b = 8'd40;  #10 
a = 8'd192; b = 8'd41;  #10 
a = 8'd192; b = 8'd42;  #10 
a = 8'd192; b = 8'd43;  #10 
a = 8'd192; b = 8'd44;  #10 
a = 8'd192; b = 8'd45;  #10 
a = 8'd192; b = 8'd46;  #10 
a = 8'd192; b = 8'd47;  #10 
a = 8'd192; b = 8'd48;  #10 
a = 8'd192; b = 8'd49;  #10 
a = 8'd192; b = 8'd50;  #10 
a = 8'd192; b = 8'd51;  #10 
a = 8'd192; b = 8'd52;  #10 
a = 8'd192; b = 8'd53;  #10 
a = 8'd192; b = 8'd54;  #10 
a = 8'd192; b = 8'd55;  #10 
a = 8'd192; b = 8'd56;  #10 
a = 8'd192; b = 8'd57;  #10 
a = 8'd192; b = 8'd58;  #10 
a = 8'd192; b = 8'd59;  #10 
a = 8'd192; b = 8'd60;  #10 
a = 8'd192; b = 8'd61;  #10 
a = 8'd192; b = 8'd62;  #10 
a = 8'd192; b = 8'd63;  #10 
a = 8'd192; b = 8'd64;  #10 
a = 8'd192; b = 8'd65;  #10 
a = 8'd192; b = 8'd66;  #10 
a = 8'd192; b = 8'd67;  #10 
a = 8'd192; b = 8'd68;  #10 
a = 8'd192; b = 8'd69;  #10 
a = 8'd192; b = 8'd70;  #10 
a = 8'd192; b = 8'd71;  #10 
a = 8'd192; b = 8'd72;  #10 
a = 8'd192; b = 8'd73;  #10 
a = 8'd192; b = 8'd74;  #10 
a = 8'd192; b = 8'd75;  #10 
a = 8'd192; b = 8'd76;  #10 
a = 8'd192; b = 8'd77;  #10 
a = 8'd192; b = 8'd78;  #10 
a = 8'd192; b = 8'd79;  #10 
a = 8'd192; b = 8'd80;  #10 
a = 8'd192; b = 8'd81;  #10 
a = 8'd192; b = 8'd82;  #10 
a = 8'd192; b = 8'd83;  #10 
a = 8'd192; b = 8'd84;  #10 
a = 8'd192; b = 8'd85;  #10 
a = 8'd192; b = 8'd86;  #10 
a = 8'd192; b = 8'd87;  #10 
a = 8'd192; b = 8'd88;  #10 
a = 8'd192; b = 8'd89;  #10 
a = 8'd192; b = 8'd90;  #10 
a = 8'd192; b = 8'd91;  #10 
a = 8'd192; b = 8'd92;  #10 
a = 8'd192; b = 8'd93;  #10 
a = 8'd192; b = 8'd94;  #10 
a = 8'd192; b = 8'd95;  #10 
a = 8'd192; b = 8'd96;  #10 
a = 8'd192; b = 8'd97;  #10 
a = 8'd192; b = 8'd98;  #10 
a = 8'd192; b = 8'd99;  #10 
a = 8'd192; b = 8'd100;  #10 
a = 8'd192; b = 8'd101;  #10 
a = 8'd192; b = 8'd102;  #10 
a = 8'd192; b = 8'd103;  #10 
a = 8'd192; b = 8'd104;  #10 
a = 8'd192; b = 8'd105;  #10 
a = 8'd192; b = 8'd106;  #10 
a = 8'd192; b = 8'd107;  #10 
a = 8'd192; b = 8'd108;  #10 
a = 8'd192; b = 8'd109;  #10 
a = 8'd192; b = 8'd110;  #10 
a = 8'd192; b = 8'd111;  #10 
a = 8'd192; b = 8'd112;  #10 
a = 8'd192; b = 8'd113;  #10 
a = 8'd192; b = 8'd114;  #10 
a = 8'd192; b = 8'd115;  #10 
a = 8'd192; b = 8'd116;  #10 
a = 8'd192; b = 8'd117;  #10 
a = 8'd192; b = 8'd118;  #10 
a = 8'd192; b = 8'd119;  #10 
a = 8'd192; b = 8'd120;  #10 
a = 8'd192; b = 8'd121;  #10 
a = 8'd192; b = 8'd122;  #10 
a = 8'd192; b = 8'd123;  #10 
a = 8'd192; b = 8'd124;  #10 
a = 8'd192; b = 8'd125;  #10 
a = 8'd192; b = 8'd126;  #10 
a = 8'd192; b = 8'd127;  #10 
a = 8'd192; b = 8'd128;  #10 
a = 8'd192; b = 8'd129;  #10 
a = 8'd192; b = 8'd130;  #10 
a = 8'd192; b = 8'd131;  #10 
a = 8'd192; b = 8'd132;  #10 
a = 8'd192; b = 8'd133;  #10 
a = 8'd192; b = 8'd134;  #10 
a = 8'd192; b = 8'd135;  #10 
a = 8'd192; b = 8'd136;  #10 
a = 8'd192; b = 8'd137;  #10 
a = 8'd192; b = 8'd138;  #10 
a = 8'd192; b = 8'd139;  #10 
a = 8'd192; b = 8'd140;  #10 
a = 8'd192; b = 8'd141;  #10 
a = 8'd192; b = 8'd142;  #10 
a = 8'd192; b = 8'd143;  #10 
a = 8'd192; b = 8'd144;  #10 
a = 8'd192; b = 8'd145;  #10 
a = 8'd192; b = 8'd146;  #10 
a = 8'd192; b = 8'd147;  #10 
a = 8'd192; b = 8'd148;  #10 
a = 8'd192; b = 8'd149;  #10 
a = 8'd192; b = 8'd150;  #10 
a = 8'd192; b = 8'd151;  #10 
a = 8'd192; b = 8'd152;  #10 
a = 8'd192; b = 8'd153;  #10 
a = 8'd192; b = 8'd154;  #10 
a = 8'd192; b = 8'd155;  #10 
a = 8'd192; b = 8'd156;  #10 
a = 8'd192; b = 8'd157;  #10 
a = 8'd192; b = 8'd158;  #10 
a = 8'd192; b = 8'd159;  #10 
a = 8'd192; b = 8'd160;  #10 
a = 8'd192; b = 8'd161;  #10 
a = 8'd192; b = 8'd162;  #10 
a = 8'd192; b = 8'd163;  #10 
a = 8'd192; b = 8'd164;  #10 
a = 8'd192; b = 8'd165;  #10 
a = 8'd192; b = 8'd166;  #10 
a = 8'd192; b = 8'd167;  #10 
a = 8'd192; b = 8'd168;  #10 
a = 8'd192; b = 8'd169;  #10 
a = 8'd192; b = 8'd170;  #10 
a = 8'd192; b = 8'd171;  #10 
a = 8'd192; b = 8'd172;  #10 
a = 8'd192; b = 8'd173;  #10 
a = 8'd192; b = 8'd174;  #10 
a = 8'd192; b = 8'd175;  #10 
a = 8'd192; b = 8'd176;  #10 
a = 8'd192; b = 8'd177;  #10 
a = 8'd192; b = 8'd178;  #10 
a = 8'd192; b = 8'd179;  #10 
a = 8'd192; b = 8'd180;  #10 
a = 8'd192; b = 8'd181;  #10 
a = 8'd192; b = 8'd182;  #10 
a = 8'd192; b = 8'd183;  #10 
a = 8'd192; b = 8'd184;  #10 
a = 8'd192; b = 8'd185;  #10 
a = 8'd192; b = 8'd186;  #10 
a = 8'd192; b = 8'd187;  #10 
a = 8'd192; b = 8'd188;  #10 
a = 8'd192; b = 8'd189;  #10 
a = 8'd192; b = 8'd190;  #10 
a = 8'd192; b = 8'd191;  #10 
a = 8'd192; b = 8'd192;  #10 
a = 8'd192; b = 8'd193;  #10 
a = 8'd192; b = 8'd194;  #10 
a = 8'd192; b = 8'd195;  #10 
a = 8'd192; b = 8'd196;  #10 
a = 8'd192; b = 8'd197;  #10 
a = 8'd192; b = 8'd198;  #10 
a = 8'd192; b = 8'd199;  #10 
a = 8'd192; b = 8'd200;  #10 
a = 8'd192; b = 8'd201;  #10 
a = 8'd192; b = 8'd202;  #10 
a = 8'd192; b = 8'd203;  #10 
a = 8'd192; b = 8'd204;  #10 
a = 8'd192; b = 8'd205;  #10 
a = 8'd192; b = 8'd206;  #10 
a = 8'd192; b = 8'd207;  #10 
a = 8'd192; b = 8'd208;  #10 
a = 8'd192; b = 8'd209;  #10 
a = 8'd192; b = 8'd210;  #10 
a = 8'd192; b = 8'd211;  #10 
a = 8'd192; b = 8'd212;  #10 
a = 8'd192; b = 8'd213;  #10 
a = 8'd192; b = 8'd214;  #10 
a = 8'd192; b = 8'd215;  #10 
a = 8'd192; b = 8'd216;  #10 
a = 8'd192; b = 8'd217;  #10 
a = 8'd192; b = 8'd218;  #10 
a = 8'd192; b = 8'd219;  #10 
a = 8'd192; b = 8'd220;  #10 
a = 8'd192; b = 8'd221;  #10 
a = 8'd192; b = 8'd222;  #10 
a = 8'd192; b = 8'd223;  #10 
a = 8'd192; b = 8'd224;  #10 
a = 8'd192; b = 8'd225;  #10 
a = 8'd192; b = 8'd226;  #10 
a = 8'd192; b = 8'd227;  #10 
a = 8'd192; b = 8'd228;  #10 
a = 8'd192; b = 8'd229;  #10 
a = 8'd192; b = 8'd230;  #10 
a = 8'd192; b = 8'd231;  #10 
a = 8'd192; b = 8'd232;  #10 
a = 8'd192; b = 8'd233;  #10 
a = 8'd192; b = 8'd234;  #10 
a = 8'd192; b = 8'd235;  #10 
a = 8'd192; b = 8'd236;  #10 
a = 8'd192; b = 8'd237;  #10 
a = 8'd192; b = 8'd238;  #10 
a = 8'd192; b = 8'd239;  #10 
a = 8'd192; b = 8'd240;  #10 
a = 8'd192; b = 8'd241;  #10 
a = 8'd192; b = 8'd242;  #10 
a = 8'd192; b = 8'd243;  #10 
a = 8'd192; b = 8'd244;  #10 
a = 8'd192; b = 8'd245;  #10 
a = 8'd192; b = 8'd246;  #10 
a = 8'd192; b = 8'd247;  #10 
a = 8'd192; b = 8'd248;  #10 
a = 8'd192; b = 8'd249;  #10 
a = 8'd192; b = 8'd250;  #10 
a = 8'd192; b = 8'd251;  #10 
a = 8'd192; b = 8'd252;  #10 
a = 8'd192; b = 8'd253;  #10 
a = 8'd192; b = 8'd254;  #10 
a = 8'd192; b = 8'd255;  #10 
a = 8'd193; b = 8'd0;  #10 
a = 8'd193; b = 8'd1;  #10 
a = 8'd193; b = 8'd2;  #10 
a = 8'd193; b = 8'd3;  #10 
a = 8'd193; b = 8'd4;  #10 
a = 8'd193; b = 8'd5;  #10 
a = 8'd193; b = 8'd6;  #10 
a = 8'd193; b = 8'd7;  #10 
a = 8'd193; b = 8'd8;  #10 
a = 8'd193; b = 8'd9;  #10 
a = 8'd193; b = 8'd10;  #10 
a = 8'd193; b = 8'd11;  #10 
a = 8'd193; b = 8'd12;  #10 
a = 8'd193; b = 8'd13;  #10 
a = 8'd193; b = 8'd14;  #10 
a = 8'd193; b = 8'd15;  #10 
a = 8'd193; b = 8'd16;  #10 
a = 8'd193; b = 8'd17;  #10 
a = 8'd193; b = 8'd18;  #10 
a = 8'd193; b = 8'd19;  #10 
a = 8'd193; b = 8'd20;  #10 
a = 8'd193; b = 8'd21;  #10 
a = 8'd193; b = 8'd22;  #10 
a = 8'd193; b = 8'd23;  #10 
a = 8'd193; b = 8'd24;  #10 
a = 8'd193; b = 8'd25;  #10 
a = 8'd193; b = 8'd26;  #10 
a = 8'd193; b = 8'd27;  #10 
a = 8'd193; b = 8'd28;  #10 
a = 8'd193; b = 8'd29;  #10 
a = 8'd193; b = 8'd30;  #10 
a = 8'd193; b = 8'd31;  #10 
a = 8'd193; b = 8'd32;  #10 
a = 8'd193; b = 8'd33;  #10 
a = 8'd193; b = 8'd34;  #10 
a = 8'd193; b = 8'd35;  #10 
a = 8'd193; b = 8'd36;  #10 
a = 8'd193; b = 8'd37;  #10 
a = 8'd193; b = 8'd38;  #10 
a = 8'd193; b = 8'd39;  #10 
a = 8'd193; b = 8'd40;  #10 
a = 8'd193; b = 8'd41;  #10 
a = 8'd193; b = 8'd42;  #10 
a = 8'd193; b = 8'd43;  #10 
a = 8'd193; b = 8'd44;  #10 
a = 8'd193; b = 8'd45;  #10 
a = 8'd193; b = 8'd46;  #10 
a = 8'd193; b = 8'd47;  #10 
a = 8'd193; b = 8'd48;  #10 
a = 8'd193; b = 8'd49;  #10 
a = 8'd193; b = 8'd50;  #10 
a = 8'd193; b = 8'd51;  #10 
a = 8'd193; b = 8'd52;  #10 
a = 8'd193; b = 8'd53;  #10 
a = 8'd193; b = 8'd54;  #10 
a = 8'd193; b = 8'd55;  #10 
a = 8'd193; b = 8'd56;  #10 
a = 8'd193; b = 8'd57;  #10 
a = 8'd193; b = 8'd58;  #10 
a = 8'd193; b = 8'd59;  #10 
a = 8'd193; b = 8'd60;  #10 
a = 8'd193; b = 8'd61;  #10 
a = 8'd193; b = 8'd62;  #10 
a = 8'd193; b = 8'd63;  #10 
a = 8'd193; b = 8'd64;  #10 
a = 8'd193; b = 8'd65;  #10 
a = 8'd193; b = 8'd66;  #10 
a = 8'd193; b = 8'd67;  #10 
a = 8'd193; b = 8'd68;  #10 
a = 8'd193; b = 8'd69;  #10 
a = 8'd193; b = 8'd70;  #10 
a = 8'd193; b = 8'd71;  #10 
a = 8'd193; b = 8'd72;  #10 
a = 8'd193; b = 8'd73;  #10 
a = 8'd193; b = 8'd74;  #10 
a = 8'd193; b = 8'd75;  #10 
a = 8'd193; b = 8'd76;  #10 
a = 8'd193; b = 8'd77;  #10 
a = 8'd193; b = 8'd78;  #10 
a = 8'd193; b = 8'd79;  #10 
a = 8'd193; b = 8'd80;  #10 
a = 8'd193; b = 8'd81;  #10 
a = 8'd193; b = 8'd82;  #10 
a = 8'd193; b = 8'd83;  #10 
a = 8'd193; b = 8'd84;  #10 
a = 8'd193; b = 8'd85;  #10 
a = 8'd193; b = 8'd86;  #10 
a = 8'd193; b = 8'd87;  #10 
a = 8'd193; b = 8'd88;  #10 
a = 8'd193; b = 8'd89;  #10 
a = 8'd193; b = 8'd90;  #10 
a = 8'd193; b = 8'd91;  #10 
a = 8'd193; b = 8'd92;  #10 
a = 8'd193; b = 8'd93;  #10 
a = 8'd193; b = 8'd94;  #10 
a = 8'd193; b = 8'd95;  #10 
a = 8'd193; b = 8'd96;  #10 
a = 8'd193; b = 8'd97;  #10 
a = 8'd193; b = 8'd98;  #10 
a = 8'd193; b = 8'd99;  #10 
a = 8'd193; b = 8'd100;  #10 
a = 8'd193; b = 8'd101;  #10 
a = 8'd193; b = 8'd102;  #10 
a = 8'd193; b = 8'd103;  #10 
a = 8'd193; b = 8'd104;  #10 
a = 8'd193; b = 8'd105;  #10 
a = 8'd193; b = 8'd106;  #10 
a = 8'd193; b = 8'd107;  #10 
a = 8'd193; b = 8'd108;  #10 
a = 8'd193; b = 8'd109;  #10 
a = 8'd193; b = 8'd110;  #10 
a = 8'd193; b = 8'd111;  #10 
a = 8'd193; b = 8'd112;  #10 
a = 8'd193; b = 8'd113;  #10 
a = 8'd193; b = 8'd114;  #10 
a = 8'd193; b = 8'd115;  #10 
a = 8'd193; b = 8'd116;  #10 
a = 8'd193; b = 8'd117;  #10 
a = 8'd193; b = 8'd118;  #10 
a = 8'd193; b = 8'd119;  #10 
a = 8'd193; b = 8'd120;  #10 
a = 8'd193; b = 8'd121;  #10 
a = 8'd193; b = 8'd122;  #10 
a = 8'd193; b = 8'd123;  #10 
a = 8'd193; b = 8'd124;  #10 
a = 8'd193; b = 8'd125;  #10 
a = 8'd193; b = 8'd126;  #10 
a = 8'd193; b = 8'd127;  #10 
a = 8'd193; b = 8'd128;  #10 
a = 8'd193; b = 8'd129;  #10 
a = 8'd193; b = 8'd130;  #10 
a = 8'd193; b = 8'd131;  #10 
a = 8'd193; b = 8'd132;  #10 
a = 8'd193; b = 8'd133;  #10 
a = 8'd193; b = 8'd134;  #10 
a = 8'd193; b = 8'd135;  #10 
a = 8'd193; b = 8'd136;  #10 
a = 8'd193; b = 8'd137;  #10 
a = 8'd193; b = 8'd138;  #10 
a = 8'd193; b = 8'd139;  #10 
a = 8'd193; b = 8'd140;  #10 
a = 8'd193; b = 8'd141;  #10 
a = 8'd193; b = 8'd142;  #10 
a = 8'd193; b = 8'd143;  #10 
a = 8'd193; b = 8'd144;  #10 
a = 8'd193; b = 8'd145;  #10 
a = 8'd193; b = 8'd146;  #10 
a = 8'd193; b = 8'd147;  #10 
a = 8'd193; b = 8'd148;  #10 
a = 8'd193; b = 8'd149;  #10 
a = 8'd193; b = 8'd150;  #10 
a = 8'd193; b = 8'd151;  #10 
a = 8'd193; b = 8'd152;  #10 
a = 8'd193; b = 8'd153;  #10 
a = 8'd193; b = 8'd154;  #10 
a = 8'd193; b = 8'd155;  #10 
a = 8'd193; b = 8'd156;  #10 
a = 8'd193; b = 8'd157;  #10 
a = 8'd193; b = 8'd158;  #10 
a = 8'd193; b = 8'd159;  #10 
a = 8'd193; b = 8'd160;  #10 
a = 8'd193; b = 8'd161;  #10 
a = 8'd193; b = 8'd162;  #10 
a = 8'd193; b = 8'd163;  #10 
a = 8'd193; b = 8'd164;  #10 
a = 8'd193; b = 8'd165;  #10 
a = 8'd193; b = 8'd166;  #10 
a = 8'd193; b = 8'd167;  #10 
a = 8'd193; b = 8'd168;  #10 
a = 8'd193; b = 8'd169;  #10 
a = 8'd193; b = 8'd170;  #10 
a = 8'd193; b = 8'd171;  #10 
a = 8'd193; b = 8'd172;  #10 
a = 8'd193; b = 8'd173;  #10 
a = 8'd193; b = 8'd174;  #10 
a = 8'd193; b = 8'd175;  #10 
a = 8'd193; b = 8'd176;  #10 
a = 8'd193; b = 8'd177;  #10 
a = 8'd193; b = 8'd178;  #10 
a = 8'd193; b = 8'd179;  #10 
a = 8'd193; b = 8'd180;  #10 
a = 8'd193; b = 8'd181;  #10 
a = 8'd193; b = 8'd182;  #10 
a = 8'd193; b = 8'd183;  #10 
a = 8'd193; b = 8'd184;  #10 
a = 8'd193; b = 8'd185;  #10 
a = 8'd193; b = 8'd186;  #10 
a = 8'd193; b = 8'd187;  #10 
a = 8'd193; b = 8'd188;  #10 
a = 8'd193; b = 8'd189;  #10 
a = 8'd193; b = 8'd190;  #10 
a = 8'd193; b = 8'd191;  #10 
a = 8'd193; b = 8'd192;  #10 
a = 8'd193; b = 8'd193;  #10 
a = 8'd193; b = 8'd194;  #10 
a = 8'd193; b = 8'd195;  #10 
a = 8'd193; b = 8'd196;  #10 
a = 8'd193; b = 8'd197;  #10 
a = 8'd193; b = 8'd198;  #10 
a = 8'd193; b = 8'd199;  #10 
a = 8'd193; b = 8'd200;  #10 
a = 8'd193; b = 8'd201;  #10 
a = 8'd193; b = 8'd202;  #10 
a = 8'd193; b = 8'd203;  #10 
a = 8'd193; b = 8'd204;  #10 
a = 8'd193; b = 8'd205;  #10 
a = 8'd193; b = 8'd206;  #10 
a = 8'd193; b = 8'd207;  #10 
a = 8'd193; b = 8'd208;  #10 
a = 8'd193; b = 8'd209;  #10 
a = 8'd193; b = 8'd210;  #10 
a = 8'd193; b = 8'd211;  #10 
a = 8'd193; b = 8'd212;  #10 
a = 8'd193; b = 8'd213;  #10 
a = 8'd193; b = 8'd214;  #10 
a = 8'd193; b = 8'd215;  #10 
a = 8'd193; b = 8'd216;  #10 
a = 8'd193; b = 8'd217;  #10 
a = 8'd193; b = 8'd218;  #10 
a = 8'd193; b = 8'd219;  #10 
a = 8'd193; b = 8'd220;  #10 
a = 8'd193; b = 8'd221;  #10 
a = 8'd193; b = 8'd222;  #10 
a = 8'd193; b = 8'd223;  #10 
a = 8'd193; b = 8'd224;  #10 
a = 8'd193; b = 8'd225;  #10 
a = 8'd193; b = 8'd226;  #10 
a = 8'd193; b = 8'd227;  #10 
a = 8'd193; b = 8'd228;  #10 
a = 8'd193; b = 8'd229;  #10 
a = 8'd193; b = 8'd230;  #10 
a = 8'd193; b = 8'd231;  #10 
a = 8'd193; b = 8'd232;  #10 
a = 8'd193; b = 8'd233;  #10 
a = 8'd193; b = 8'd234;  #10 
a = 8'd193; b = 8'd235;  #10 
a = 8'd193; b = 8'd236;  #10 
a = 8'd193; b = 8'd237;  #10 
a = 8'd193; b = 8'd238;  #10 
a = 8'd193; b = 8'd239;  #10 
a = 8'd193; b = 8'd240;  #10 
a = 8'd193; b = 8'd241;  #10 
a = 8'd193; b = 8'd242;  #10 
a = 8'd193; b = 8'd243;  #10 
a = 8'd193; b = 8'd244;  #10 
a = 8'd193; b = 8'd245;  #10 
a = 8'd193; b = 8'd246;  #10 
a = 8'd193; b = 8'd247;  #10 
a = 8'd193; b = 8'd248;  #10 
a = 8'd193; b = 8'd249;  #10 
a = 8'd193; b = 8'd250;  #10 
a = 8'd193; b = 8'd251;  #10 
a = 8'd193; b = 8'd252;  #10 
a = 8'd193; b = 8'd253;  #10 
a = 8'd193; b = 8'd254;  #10 
a = 8'd193; b = 8'd255;  #10 
a = 8'd194; b = 8'd0;  #10 
a = 8'd194; b = 8'd1;  #10 
a = 8'd194; b = 8'd2;  #10 
a = 8'd194; b = 8'd3;  #10 
a = 8'd194; b = 8'd4;  #10 
a = 8'd194; b = 8'd5;  #10 
a = 8'd194; b = 8'd6;  #10 
a = 8'd194; b = 8'd7;  #10 
a = 8'd194; b = 8'd8;  #10 
a = 8'd194; b = 8'd9;  #10 
a = 8'd194; b = 8'd10;  #10 
a = 8'd194; b = 8'd11;  #10 
a = 8'd194; b = 8'd12;  #10 
a = 8'd194; b = 8'd13;  #10 
a = 8'd194; b = 8'd14;  #10 
a = 8'd194; b = 8'd15;  #10 
a = 8'd194; b = 8'd16;  #10 
a = 8'd194; b = 8'd17;  #10 
a = 8'd194; b = 8'd18;  #10 
a = 8'd194; b = 8'd19;  #10 
a = 8'd194; b = 8'd20;  #10 
a = 8'd194; b = 8'd21;  #10 
a = 8'd194; b = 8'd22;  #10 
a = 8'd194; b = 8'd23;  #10 
a = 8'd194; b = 8'd24;  #10 
a = 8'd194; b = 8'd25;  #10 
a = 8'd194; b = 8'd26;  #10 
a = 8'd194; b = 8'd27;  #10 
a = 8'd194; b = 8'd28;  #10 
a = 8'd194; b = 8'd29;  #10 
a = 8'd194; b = 8'd30;  #10 
a = 8'd194; b = 8'd31;  #10 
a = 8'd194; b = 8'd32;  #10 
a = 8'd194; b = 8'd33;  #10 
a = 8'd194; b = 8'd34;  #10 
a = 8'd194; b = 8'd35;  #10 
a = 8'd194; b = 8'd36;  #10 
a = 8'd194; b = 8'd37;  #10 
a = 8'd194; b = 8'd38;  #10 
a = 8'd194; b = 8'd39;  #10 
a = 8'd194; b = 8'd40;  #10 
a = 8'd194; b = 8'd41;  #10 
a = 8'd194; b = 8'd42;  #10 
a = 8'd194; b = 8'd43;  #10 
a = 8'd194; b = 8'd44;  #10 
a = 8'd194; b = 8'd45;  #10 
a = 8'd194; b = 8'd46;  #10 
a = 8'd194; b = 8'd47;  #10 
a = 8'd194; b = 8'd48;  #10 
a = 8'd194; b = 8'd49;  #10 
a = 8'd194; b = 8'd50;  #10 
a = 8'd194; b = 8'd51;  #10 
a = 8'd194; b = 8'd52;  #10 
a = 8'd194; b = 8'd53;  #10 
a = 8'd194; b = 8'd54;  #10 
a = 8'd194; b = 8'd55;  #10 
a = 8'd194; b = 8'd56;  #10 
a = 8'd194; b = 8'd57;  #10 
a = 8'd194; b = 8'd58;  #10 
a = 8'd194; b = 8'd59;  #10 
a = 8'd194; b = 8'd60;  #10 
a = 8'd194; b = 8'd61;  #10 
a = 8'd194; b = 8'd62;  #10 
a = 8'd194; b = 8'd63;  #10 
a = 8'd194; b = 8'd64;  #10 
a = 8'd194; b = 8'd65;  #10 
a = 8'd194; b = 8'd66;  #10 
a = 8'd194; b = 8'd67;  #10 
a = 8'd194; b = 8'd68;  #10 
a = 8'd194; b = 8'd69;  #10 
a = 8'd194; b = 8'd70;  #10 
a = 8'd194; b = 8'd71;  #10 
a = 8'd194; b = 8'd72;  #10 
a = 8'd194; b = 8'd73;  #10 
a = 8'd194; b = 8'd74;  #10 
a = 8'd194; b = 8'd75;  #10 
a = 8'd194; b = 8'd76;  #10 
a = 8'd194; b = 8'd77;  #10 
a = 8'd194; b = 8'd78;  #10 
a = 8'd194; b = 8'd79;  #10 
a = 8'd194; b = 8'd80;  #10 
a = 8'd194; b = 8'd81;  #10 
a = 8'd194; b = 8'd82;  #10 
a = 8'd194; b = 8'd83;  #10 
a = 8'd194; b = 8'd84;  #10 
a = 8'd194; b = 8'd85;  #10 
a = 8'd194; b = 8'd86;  #10 
a = 8'd194; b = 8'd87;  #10 
a = 8'd194; b = 8'd88;  #10 
a = 8'd194; b = 8'd89;  #10 
a = 8'd194; b = 8'd90;  #10 
a = 8'd194; b = 8'd91;  #10 
a = 8'd194; b = 8'd92;  #10 
a = 8'd194; b = 8'd93;  #10 
a = 8'd194; b = 8'd94;  #10 
a = 8'd194; b = 8'd95;  #10 
a = 8'd194; b = 8'd96;  #10 
a = 8'd194; b = 8'd97;  #10 
a = 8'd194; b = 8'd98;  #10 
a = 8'd194; b = 8'd99;  #10 
a = 8'd194; b = 8'd100;  #10 
a = 8'd194; b = 8'd101;  #10 
a = 8'd194; b = 8'd102;  #10 
a = 8'd194; b = 8'd103;  #10 
a = 8'd194; b = 8'd104;  #10 
a = 8'd194; b = 8'd105;  #10 
a = 8'd194; b = 8'd106;  #10 
a = 8'd194; b = 8'd107;  #10 
a = 8'd194; b = 8'd108;  #10 
a = 8'd194; b = 8'd109;  #10 
a = 8'd194; b = 8'd110;  #10 
a = 8'd194; b = 8'd111;  #10 
a = 8'd194; b = 8'd112;  #10 
a = 8'd194; b = 8'd113;  #10 
a = 8'd194; b = 8'd114;  #10 
a = 8'd194; b = 8'd115;  #10 
a = 8'd194; b = 8'd116;  #10 
a = 8'd194; b = 8'd117;  #10 
a = 8'd194; b = 8'd118;  #10 
a = 8'd194; b = 8'd119;  #10 
a = 8'd194; b = 8'd120;  #10 
a = 8'd194; b = 8'd121;  #10 
a = 8'd194; b = 8'd122;  #10 
a = 8'd194; b = 8'd123;  #10 
a = 8'd194; b = 8'd124;  #10 
a = 8'd194; b = 8'd125;  #10 
a = 8'd194; b = 8'd126;  #10 
a = 8'd194; b = 8'd127;  #10 
a = 8'd194; b = 8'd128;  #10 
a = 8'd194; b = 8'd129;  #10 
a = 8'd194; b = 8'd130;  #10 
a = 8'd194; b = 8'd131;  #10 
a = 8'd194; b = 8'd132;  #10 
a = 8'd194; b = 8'd133;  #10 
a = 8'd194; b = 8'd134;  #10 
a = 8'd194; b = 8'd135;  #10 
a = 8'd194; b = 8'd136;  #10 
a = 8'd194; b = 8'd137;  #10 
a = 8'd194; b = 8'd138;  #10 
a = 8'd194; b = 8'd139;  #10 
a = 8'd194; b = 8'd140;  #10 
a = 8'd194; b = 8'd141;  #10 
a = 8'd194; b = 8'd142;  #10 
a = 8'd194; b = 8'd143;  #10 
a = 8'd194; b = 8'd144;  #10 
a = 8'd194; b = 8'd145;  #10 
a = 8'd194; b = 8'd146;  #10 
a = 8'd194; b = 8'd147;  #10 
a = 8'd194; b = 8'd148;  #10 
a = 8'd194; b = 8'd149;  #10 
a = 8'd194; b = 8'd150;  #10 
a = 8'd194; b = 8'd151;  #10 
a = 8'd194; b = 8'd152;  #10 
a = 8'd194; b = 8'd153;  #10 
a = 8'd194; b = 8'd154;  #10 
a = 8'd194; b = 8'd155;  #10 
a = 8'd194; b = 8'd156;  #10 
a = 8'd194; b = 8'd157;  #10 
a = 8'd194; b = 8'd158;  #10 
a = 8'd194; b = 8'd159;  #10 
a = 8'd194; b = 8'd160;  #10 
a = 8'd194; b = 8'd161;  #10 
a = 8'd194; b = 8'd162;  #10 
a = 8'd194; b = 8'd163;  #10 
a = 8'd194; b = 8'd164;  #10 
a = 8'd194; b = 8'd165;  #10 
a = 8'd194; b = 8'd166;  #10 
a = 8'd194; b = 8'd167;  #10 
a = 8'd194; b = 8'd168;  #10 
a = 8'd194; b = 8'd169;  #10 
a = 8'd194; b = 8'd170;  #10 
a = 8'd194; b = 8'd171;  #10 
a = 8'd194; b = 8'd172;  #10 
a = 8'd194; b = 8'd173;  #10 
a = 8'd194; b = 8'd174;  #10 
a = 8'd194; b = 8'd175;  #10 
a = 8'd194; b = 8'd176;  #10 
a = 8'd194; b = 8'd177;  #10 
a = 8'd194; b = 8'd178;  #10 
a = 8'd194; b = 8'd179;  #10 
a = 8'd194; b = 8'd180;  #10 
a = 8'd194; b = 8'd181;  #10 
a = 8'd194; b = 8'd182;  #10 
a = 8'd194; b = 8'd183;  #10 
a = 8'd194; b = 8'd184;  #10 
a = 8'd194; b = 8'd185;  #10 
a = 8'd194; b = 8'd186;  #10 
a = 8'd194; b = 8'd187;  #10 
a = 8'd194; b = 8'd188;  #10 
a = 8'd194; b = 8'd189;  #10 
a = 8'd194; b = 8'd190;  #10 
a = 8'd194; b = 8'd191;  #10 
a = 8'd194; b = 8'd192;  #10 
a = 8'd194; b = 8'd193;  #10 
a = 8'd194; b = 8'd194;  #10 
a = 8'd194; b = 8'd195;  #10 
a = 8'd194; b = 8'd196;  #10 
a = 8'd194; b = 8'd197;  #10 
a = 8'd194; b = 8'd198;  #10 
a = 8'd194; b = 8'd199;  #10 
a = 8'd194; b = 8'd200;  #10 
a = 8'd194; b = 8'd201;  #10 
a = 8'd194; b = 8'd202;  #10 
a = 8'd194; b = 8'd203;  #10 
a = 8'd194; b = 8'd204;  #10 
a = 8'd194; b = 8'd205;  #10 
a = 8'd194; b = 8'd206;  #10 
a = 8'd194; b = 8'd207;  #10 
a = 8'd194; b = 8'd208;  #10 
a = 8'd194; b = 8'd209;  #10 
a = 8'd194; b = 8'd210;  #10 
a = 8'd194; b = 8'd211;  #10 
a = 8'd194; b = 8'd212;  #10 
a = 8'd194; b = 8'd213;  #10 
a = 8'd194; b = 8'd214;  #10 
a = 8'd194; b = 8'd215;  #10 
a = 8'd194; b = 8'd216;  #10 
a = 8'd194; b = 8'd217;  #10 
a = 8'd194; b = 8'd218;  #10 
a = 8'd194; b = 8'd219;  #10 
a = 8'd194; b = 8'd220;  #10 
a = 8'd194; b = 8'd221;  #10 
a = 8'd194; b = 8'd222;  #10 
a = 8'd194; b = 8'd223;  #10 
a = 8'd194; b = 8'd224;  #10 
a = 8'd194; b = 8'd225;  #10 
a = 8'd194; b = 8'd226;  #10 
a = 8'd194; b = 8'd227;  #10 
a = 8'd194; b = 8'd228;  #10 
a = 8'd194; b = 8'd229;  #10 
a = 8'd194; b = 8'd230;  #10 
a = 8'd194; b = 8'd231;  #10 
a = 8'd194; b = 8'd232;  #10 
a = 8'd194; b = 8'd233;  #10 
a = 8'd194; b = 8'd234;  #10 
a = 8'd194; b = 8'd235;  #10 
a = 8'd194; b = 8'd236;  #10 
a = 8'd194; b = 8'd237;  #10 
a = 8'd194; b = 8'd238;  #10 
a = 8'd194; b = 8'd239;  #10 
a = 8'd194; b = 8'd240;  #10 
a = 8'd194; b = 8'd241;  #10 
a = 8'd194; b = 8'd242;  #10 
a = 8'd194; b = 8'd243;  #10 
a = 8'd194; b = 8'd244;  #10 
a = 8'd194; b = 8'd245;  #10 
a = 8'd194; b = 8'd246;  #10 
a = 8'd194; b = 8'd247;  #10 
a = 8'd194; b = 8'd248;  #10 
a = 8'd194; b = 8'd249;  #10 
a = 8'd194; b = 8'd250;  #10 
a = 8'd194; b = 8'd251;  #10 
a = 8'd194; b = 8'd252;  #10 
a = 8'd194; b = 8'd253;  #10 
a = 8'd194; b = 8'd254;  #10 
a = 8'd194; b = 8'd255;  #10 
a = 8'd195; b = 8'd0;  #10 
a = 8'd195; b = 8'd1;  #10 
a = 8'd195; b = 8'd2;  #10 
a = 8'd195; b = 8'd3;  #10 
a = 8'd195; b = 8'd4;  #10 
a = 8'd195; b = 8'd5;  #10 
a = 8'd195; b = 8'd6;  #10 
a = 8'd195; b = 8'd7;  #10 
a = 8'd195; b = 8'd8;  #10 
a = 8'd195; b = 8'd9;  #10 
a = 8'd195; b = 8'd10;  #10 
a = 8'd195; b = 8'd11;  #10 
a = 8'd195; b = 8'd12;  #10 
a = 8'd195; b = 8'd13;  #10 
a = 8'd195; b = 8'd14;  #10 
a = 8'd195; b = 8'd15;  #10 
a = 8'd195; b = 8'd16;  #10 
a = 8'd195; b = 8'd17;  #10 
a = 8'd195; b = 8'd18;  #10 
a = 8'd195; b = 8'd19;  #10 
a = 8'd195; b = 8'd20;  #10 
a = 8'd195; b = 8'd21;  #10 
a = 8'd195; b = 8'd22;  #10 
a = 8'd195; b = 8'd23;  #10 
a = 8'd195; b = 8'd24;  #10 
a = 8'd195; b = 8'd25;  #10 
a = 8'd195; b = 8'd26;  #10 
a = 8'd195; b = 8'd27;  #10 
a = 8'd195; b = 8'd28;  #10 
a = 8'd195; b = 8'd29;  #10 
a = 8'd195; b = 8'd30;  #10 
a = 8'd195; b = 8'd31;  #10 
a = 8'd195; b = 8'd32;  #10 
a = 8'd195; b = 8'd33;  #10 
a = 8'd195; b = 8'd34;  #10 
a = 8'd195; b = 8'd35;  #10 
a = 8'd195; b = 8'd36;  #10 
a = 8'd195; b = 8'd37;  #10 
a = 8'd195; b = 8'd38;  #10 
a = 8'd195; b = 8'd39;  #10 
a = 8'd195; b = 8'd40;  #10 
a = 8'd195; b = 8'd41;  #10 
a = 8'd195; b = 8'd42;  #10 
a = 8'd195; b = 8'd43;  #10 
a = 8'd195; b = 8'd44;  #10 
a = 8'd195; b = 8'd45;  #10 
a = 8'd195; b = 8'd46;  #10 
a = 8'd195; b = 8'd47;  #10 
a = 8'd195; b = 8'd48;  #10 
a = 8'd195; b = 8'd49;  #10 
a = 8'd195; b = 8'd50;  #10 
a = 8'd195; b = 8'd51;  #10 
a = 8'd195; b = 8'd52;  #10 
a = 8'd195; b = 8'd53;  #10 
a = 8'd195; b = 8'd54;  #10 
a = 8'd195; b = 8'd55;  #10 
a = 8'd195; b = 8'd56;  #10 
a = 8'd195; b = 8'd57;  #10 
a = 8'd195; b = 8'd58;  #10 
a = 8'd195; b = 8'd59;  #10 
a = 8'd195; b = 8'd60;  #10 
a = 8'd195; b = 8'd61;  #10 
a = 8'd195; b = 8'd62;  #10 
a = 8'd195; b = 8'd63;  #10 
a = 8'd195; b = 8'd64;  #10 
a = 8'd195; b = 8'd65;  #10 
a = 8'd195; b = 8'd66;  #10 
a = 8'd195; b = 8'd67;  #10 
a = 8'd195; b = 8'd68;  #10 
a = 8'd195; b = 8'd69;  #10 
a = 8'd195; b = 8'd70;  #10 
a = 8'd195; b = 8'd71;  #10 
a = 8'd195; b = 8'd72;  #10 
a = 8'd195; b = 8'd73;  #10 
a = 8'd195; b = 8'd74;  #10 
a = 8'd195; b = 8'd75;  #10 
a = 8'd195; b = 8'd76;  #10 
a = 8'd195; b = 8'd77;  #10 
a = 8'd195; b = 8'd78;  #10 
a = 8'd195; b = 8'd79;  #10 
a = 8'd195; b = 8'd80;  #10 
a = 8'd195; b = 8'd81;  #10 
a = 8'd195; b = 8'd82;  #10 
a = 8'd195; b = 8'd83;  #10 
a = 8'd195; b = 8'd84;  #10 
a = 8'd195; b = 8'd85;  #10 
a = 8'd195; b = 8'd86;  #10 
a = 8'd195; b = 8'd87;  #10 
a = 8'd195; b = 8'd88;  #10 
a = 8'd195; b = 8'd89;  #10 
a = 8'd195; b = 8'd90;  #10 
a = 8'd195; b = 8'd91;  #10 
a = 8'd195; b = 8'd92;  #10 
a = 8'd195; b = 8'd93;  #10 
a = 8'd195; b = 8'd94;  #10 
a = 8'd195; b = 8'd95;  #10 
a = 8'd195; b = 8'd96;  #10 
a = 8'd195; b = 8'd97;  #10 
a = 8'd195; b = 8'd98;  #10 
a = 8'd195; b = 8'd99;  #10 
a = 8'd195; b = 8'd100;  #10 
a = 8'd195; b = 8'd101;  #10 
a = 8'd195; b = 8'd102;  #10 
a = 8'd195; b = 8'd103;  #10 
a = 8'd195; b = 8'd104;  #10 
a = 8'd195; b = 8'd105;  #10 
a = 8'd195; b = 8'd106;  #10 
a = 8'd195; b = 8'd107;  #10 
a = 8'd195; b = 8'd108;  #10 
a = 8'd195; b = 8'd109;  #10 
a = 8'd195; b = 8'd110;  #10 
a = 8'd195; b = 8'd111;  #10 
a = 8'd195; b = 8'd112;  #10 
a = 8'd195; b = 8'd113;  #10 
a = 8'd195; b = 8'd114;  #10 
a = 8'd195; b = 8'd115;  #10 
a = 8'd195; b = 8'd116;  #10 
a = 8'd195; b = 8'd117;  #10 
a = 8'd195; b = 8'd118;  #10 
a = 8'd195; b = 8'd119;  #10 
a = 8'd195; b = 8'd120;  #10 
a = 8'd195; b = 8'd121;  #10 
a = 8'd195; b = 8'd122;  #10 
a = 8'd195; b = 8'd123;  #10 
a = 8'd195; b = 8'd124;  #10 
a = 8'd195; b = 8'd125;  #10 
a = 8'd195; b = 8'd126;  #10 
a = 8'd195; b = 8'd127;  #10 
a = 8'd195; b = 8'd128;  #10 
a = 8'd195; b = 8'd129;  #10 
a = 8'd195; b = 8'd130;  #10 
a = 8'd195; b = 8'd131;  #10 
a = 8'd195; b = 8'd132;  #10 
a = 8'd195; b = 8'd133;  #10 
a = 8'd195; b = 8'd134;  #10 
a = 8'd195; b = 8'd135;  #10 
a = 8'd195; b = 8'd136;  #10 
a = 8'd195; b = 8'd137;  #10 
a = 8'd195; b = 8'd138;  #10 
a = 8'd195; b = 8'd139;  #10 
a = 8'd195; b = 8'd140;  #10 
a = 8'd195; b = 8'd141;  #10 
a = 8'd195; b = 8'd142;  #10 
a = 8'd195; b = 8'd143;  #10 
a = 8'd195; b = 8'd144;  #10 
a = 8'd195; b = 8'd145;  #10 
a = 8'd195; b = 8'd146;  #10 
a = 8'd195; b = 8'd147;  #10 
a = 8'd195; b = 8'd148;  #10 
a = 8'd195; b = 8'd149;  #10 
a = 8'd195; b = 8'd150;  #10 
a = 8'd195; b = 8'd151;  #10 
a = 8'd195; b = 8'd152;  #10 
a = 8'd195; b = 8'd153;  #10 
a = 8'd195; b = 8'd154;  #10 
a = 8'd195; b = 8'd155;  #10 
a = 8'd195; b = 8'd156;  #10 
a = 8'd195; b = 8'd157;  #10 
a = 8'd195; b = 8'd158;  #10 
a = 8'd195; b = 8'd159;  #10 
a = 8'd195; b = 8'd160;  #10 
a = 8'd195; b = 8'd161;  #10 
a = 8'd195; b = 8'd162;  #10 
a = 8'd195; b = 8'd163;  #10 
a = 8'd195; b = 8'd164;  #10 
a = 8'd195; b = 8'd165;  #10 
a = 8'd195; b = 8'd166;  #10 
a = 8'd195; b = 8'd167;  #10 
a = 8'd195; b = 8'd168;  #10 
a = 8'd195; b = 8'd169;  #10 
a = 8'd195; b = 8'd170;  #10 
a = 8'd195; b = 8'd171;  #10 
a = 8'd195; b = 8'd172;  #10 
a = 8'd195; b = 8'd173;  #10 
a = 8'd195; b = 8'd174;  #10 
a = 8'd195; b = 8'd175;  #10 
a = 8'd195; b = 8'd176;  #10 
a = 8'd195; b = 8'd177;  #10 
a = 8'd195; b = 8'd178;  #10 
a = 8'd195; b = 8'd179;  #10 
a = 8'd195; b = 8'd180;  #10 
a = 8'd195; b = 8'd181;  #10 
a = 8'd195; b = 8'd182;  #10 
a = 8'd195; b = 8'd183;  #10 
a = 8'd195; b = 8'd184;  #10 
a = 8'd195; b = 8'd185;  #10 
a = 8'd195; b = 8'd186;  #10 
a = 8'd195; b = 8'd187;  #10 
a = 8'd195; b = 8'd188;  #10 
a = 8'd195; b = 8'd189;  #10 
a = 8'd195; b = 8'd190;  #10 
a = 8'd195; b = 8'd191;  #10 
a = 8'd195; b = 8'd192;  #10 
a = 8'd195; b = 8'd193;  #10 
a = 8'd195; b = 8'd194;  #10 
a = 8'd195; b = 8'd195;  #10 
a = 8'd195; b = 8'd196;  #10 
a = 8'd195; b = 8'd197;  #10 
a = 8'd195; b = 8'd198;  #10 
a = 8'd195; b = 8'd199;  #10 
a = 8'd195; b = 8'd200;  #10 
a = 8'd195; b = 8'd201;  #10 
a = 8'd195; b = 8'd202;  #10 
a = 8'd195; b = 8'd203;  #10 
a = 8'd195; b = 8'd204;  #10 
a = 8'd195; b = 8'd205;  #10 
a = 8'd195; b = 8'd206;  #10 
a = 8'd195; b = 8'd207;  #10 
a = 8'd195; b = 8'd208;  #10 
a = 8'd195; b = 8'd209;  #10 
a = 8'd195; b = 8'd210;  #10 
a = 8'd195; b = 8'd211;  #10 
a = 8'd195; b = 8'd212;  #10 
a = 8'd195; b = 8'd213;  #10 
a = 8'd195; b = 8'd214;  #10 
a = 8'd195; b = 8'd215;  #10 
a = 8'd195; b = 8'd216;  #10 
a = 8'd195; b = 8'd217;  #10 
a = 8'd195; b = 8'd218;  #10 
a = 8'd195; b = 8'd219;  #10 
a = 8'd195; b = 8'd220;  #10 
a = 8'd195; b = 8'd221;  #10 
a = 8'd195; b = 8'd222;  #10 
a = 8'd195; b = 8'd223;  #10 
a = 8'd195; b = 8'd224;  #10 
a = 8'd195; b = 8'd225;  #10 
a = 8'd195; b = 8'd226;  #10 
a = 8'd195; b = 8'd227;  #10 
a = 8'd195; b = 8'd228;  #10 
a = 8'd195; b = 8'd229;  #10 
a = 8'd195; b = 8'd230;  #10 
a = 8'd195; b = 8'd231;  #10 
a = 8'd195; b = 8'd232;  #10 
a = 8'd195; b = 8'd233;  #10 
a = 8'd195; b = 8'd234;  #10 
a = 8'd195; b = 8'd235;  #10 
a = 8'd195; b = 8'd236;  #10 
a = 8'd195; b = 8'd237;  #10 
a = 8'd195; b = 8'd238;  #10 
a = 8'd195; b = 8'd239;  #10 
a = 8'd195; b = 8'd240;  #10 
a = 8'd195; b = 8'd241;  #10 
a = 8'd195; b = 8'd242;  #10 
a = 8'd195; b = 8'd243;  #10 
a = 8'd195; b = 8'd244;  #10 
a = 8'd195; b = 8'd245;  #10 
a = 8'd195; b = 8'd246;  #10 
a = 8'd195; b = 8'd247;  #10 
a = 8'd195; b = 8'd248;  #10 
a = 8'd195; b = 8'd249;  #10 
a = 8'd195; b = 8'd250;  #10 
a = 8'd195; b = 8'd251;  #10 
a = 8'd195; b = 8'd252;  #10 
a = 8'd195; b = 8'd253;  #10 
a = 8'd195; b = 8'd254;  #10 
a = 8'd195; b = 8'd255;  #10 
a = 8'd196; b = 8'd0;  #10 
a = 8'd196; b = 8'd1;  #10 
a = 8'd196; b = 8'd2;  #10 
a = 8'd196; b = 8'd3;  #10 
a = 8'd196; b = 8'd4;  #10 
a = 8'd196; b = 8'd5;  #10 
a = 8'd196; b = 8'd6;  #10 
a = 8'd196; b = 8'd7;  #10 
a = 8'd196; b = 8'd8;  #10 
a = 8'd196; b = 8'd9;  #10 
a = 8'd196; b = 8'd10;  #10 
a = 8'd196; b = 8'd11;  #10 
a = 8'd196; b = 8'd12;  #10 
a = 8'd196; b = 8'd13;  #10 
a = 8'd196; b = 8'd14;  #10 
a = 8'd196; b = 8'd15;  #10 
a = 8'd196; b = 8'd16;  #10 
a = 8'd196; b = 8'd17;  #10 
a = 8'd196; b = 8'd18;  #10 
a = 8'd196; b = 8'd19;  #10 
a = 8'd196; b = 8'd20;  #10 
a = 8'd196; b = 8'd21;  #10 
a = 8'd196; b = 8'd22;  #10 
a = 8'd196; b = 8'd23;  #10 
a = 8'd196; b = 8'd24;  #10 
a = 8'd196; b = 8'd25;  #10 
a = 8'd196; b = 8'd26;  #10 
a = 8'd196; b = 8'd27;  #10 
a = 8'd196; b = 8'd28;  #10 
a = 8'd196; b = 8'd29;  #10 
a = 8'd196; b = 8'd30;  #10 
a = 8'd196; b = 8'd31;  #10 
a = 8'd196; b = 8'd32;  #10 
a = 8'd196; b = 8'd33;  #10 
a = 8'd196; b = 8'd34;  #10 
a = 8'd196; b = 8'd35;  #10 
a = 8'd196; b = 8'd36;  #10 
a = 8'd196; b = 8'd37;  #10 
a = 8'd196; b = 8'd38;  #10 
a = 8'd196; b = 8'd39;  #10 
a = 8'd196; b = 8'd40;  #10 
a = 8'd196; b = 8'd41;  #10 
a = 8'd196; b = 8'd42;  #10 
a = 8'd196; b = 8'd43;  #10 
a = 8'd196; b = 8'd44;  #10 
a = 8'd196; b = 8'd45;  #10 
a = 8'd196; b = 8'd46;  #10 
a = 8'd196; b = 8'd47;  #10 
a = 8'd196; b = 8'd48;  #10 
a = 8'd196; b = 8'd49;  #10 
a = 8'd196; b = 8'd50;  #10 
a = 8'd196; b = 8'd51;  #10 
a = 8'd196; b = 8'd52;  #10 
a = 8'd196; b = 8'd53;  #10 
a = 8'd196; b = 8'd54;  #10 
a = 8'd196; b = 8'd55;  #10 
a = 8'd196; b = 8'd56;  #10 
a = 8'd196; b = 8'd57;  #10 
a = 8'd196; b = 8'd58;  #10 
a = 8'd196; b = 8'd59;  #10 
a = 8'd196; b = 8'd60;  #10 
a = 8'd196; b = 8'd61;  #10 
a = 8'd196; b = 8'd62;  #10 
a = 8'd196; b = 8'd63;  #10 
a = 8'd196; b = 8'd64;  #10 
a = 8'd196; b = 8'd65;  #10 
a = 8'd196; b = 8'd66;  #10 
a = 8'd196; b = 8'd67;  #10 
a = 8'd196; b = 8'd68;  #10 
a = 8'd196; b = 8'd69;  #10 
a = 8'd196; b = 8'd70;  #10 
a = 8'd196; b = 8'd71;  #10 
a = 8'd196; b = 8'd72;  #10 
a = 8'd196; b = 8'd73;  #10 
a = 8'd196; b = 8'd74;  #10 
a = 8'd196; b = 8'd75;  #10 
a = 8'd196; b = 8'd76;  #10 
a = 8'd196; b = 8'd77;  #10 
a = 8'd196; b = 8'd78;  #10 
a = 8'd196; b = 8'd79;  #10 
a = 8'd196; b = 8'd80;  #10 
a = 8'd196; b = 8'd81;  #10 
a = 8'd196; b = 8'd82;  #10 
a = 8'd196; b = 8'd83;  #10 
a = 8'd196; b = 8'd84;  #10 
a = 8'd196; b = 8'd85;  #10 
a = 8'd196; b = 8'd86;  #10 
a = 8'd196; b = 8'd87;  #10 
a = 8'd196; b = 8'd88;  #10 
a = 8'd196; b = 8'd89;  #10 
a = 8'd196; b = 8'd90;  #10 
a = 8'd196; b = 8'd91;  #10 
a = 8'd196; b = 8'd92;  #10 
a = 8'd196; b = 8'd93;  #10 
a = 8'd196; b = 8'd94;  #10 
a = 8'd196; b = 8'd95;  #10 
a = 8'd196; b = 8'd96;  #10 
a = 8'd196; b = 8'd97;  #10 
a = 8'd196; b = 8'd98;  #10 
a = 8'd196; b = 8'd99;  #10 
a = 8'd196; b = 8'd100;  #10 
a = 8'd196; b = 8'd101;  #10 
a = 8'd196; b = 8'd102;  #10 
a = 8'd196; b = 8'd103;  #10 
a = 8'd196; b = 8'd104;  #10 
a = 8'd196; b = 8'd105;  #10 
a = 8'd196; b = 8'd106;  #10 
a = 8'd196; b = 8'd107;  #10 
a = 8'd196; b = 8'd108;  #10 
a = 8'd196; b = 8'd109;  #10 
a = 8'd196; b = 8'd110;  #10 
a = 8'd196; b = 8'd111;  #10 
a = 8'd196; b = 8'd112;  #10 
a = 8'd196; b = 8'd113;  #10 
a = 8'd196; b = 8'd114;  #10 
a = 8'd196; b = 8'd115;  #10 
a = 8'd196; b = 8'd116;  #10 
a = 8'd196; b = 8'd117;  #10 
a = 8'd196; b = 8'd118;  #10 
a = 8'd196; b = 8'd119;  #10 
a = 8'd196; b = 8'd120;  #10 
a = 8'd196; b = 8'd121;  #10 
a = 8'd196; b = 8'd122;  #10 
a = 8'd196; b = 8'd123;  #10 
a = 8'd196; b = 8'd124;  #10 
a = 8'd196; b = 8'd125;  #10 
a = 8'd196; b = 8'd126;  #10 
a = 8'd196; b = 8'd127;  #10 
a = 8'd196; b = 8'd128;  #10 
a = 8'd196; b = 8'd129;  #10 
a = 8'd196; b = 8'd130;  #10 
a = 8'd196; b = 8'd131;  #10 
a = 8'd196; b = 8'd132;  #10 
a = 8'd196; b = 8'd133;  #10 
a = 8'd196; b = 8'd134;  #10 
a = 8'd196; b = 8'd135;  #10 
a = 8'd196; b = 8'd136;  #10 
a = 8'd196; b = 8'd137;  #10 
a = 8'd196; b = 8'd138;  #10 
a = 8'd196; b = 8'd139;  #10 
a = 8'd196; b = 8'd140;  #10 
a = 8'd196; b = 8'd141;  #10 
a = 8'd196; b = 8'd142;  #10 
a = 8'd196; b = 8'd143;  #10 
a = 8'd196; b = 8'd144;  #10 
a = 8'd196; b = 8'd145;  #10 
a = 8'd196; b = 8'd146;  #10 
a = 8'd196; b = 8'd147;  #10 
a = 8'd196; b = 8'd148;  #10 
a = 8'd196; b = 8'd149;  #10 
a = 8'd196; b = 8'd150;  #10 
a = 8'd196; b = 8'd151;  #10 
a = 8'd196; b = 8'd152;  #10 
a = 8'd196; b = 8'd153;  #10 
a = 8'd196; b = 8'd154;  #10 
a = 8'd196; b = 8'd155;  #10 
a = 8'd196; b = 8'd156;  #10 
a = 8'd196; b = 8'd157;  #10 
a = 8'd196; b = 8'd158;  #10 
a = 8'd196; b = 8'd159;  #10 
a = 8'd196; b = 8'd160;  #10 
a = 8'd196; b = 8'd161;  #10 
a = 8'd196; b = 8'd162;  #10 
a = 8'd196; b = 8'd163;  #10 
a = 8'd196; b = 8'd164;  #10 
a = 8'd196; b = 8'd165;  #10 
a = 8'd196; b = 8'd166;  #10 
a = 8'd196; b = 8'd167;  #10 
a = 8'd196; b = 8'd168;  #10 
a = 8'd196; b = 8'd169;  #10 
a = 8'd196; b = 8'd170;  #10 
a = 8'd196; b = 8'd171;  #10 
a = 8'd196; b = 8'd172;  #10 
a = 8'd196; b = 8'd173;  #10 
a = 8'd196; b = 8'd174;  #10 
a = 8'd196; b = 8'd175;  #10 
a = 8'd196; b = 8'd176;  #10 
a = 8'd196; b = 8'd177;  #10 
a = 8'd196; b = 8'd178;  #10 
a = 8'd196; b = 8'd179;  #10 
a = 8'd196; b = 8'd180;  #10 
a = 8'd196; b = 8'd181;  #10 
a = 8'd196; b = 8'd182;  #10 
a = 8'd196; b = 8'd183;  #10 
a = 8'd196; b = 8'd184;  #10 
a = 8'd196; b = 8'd185;  #10 
a = 8'd196; b = 8'd186;  #10 
a = 8'd196; b = 8'd187;  #10 
a = 8'd196; b = 8'd188;  #10 
a = 8'd196; b = 8'd189;  #10 
a = 8'd196; b = 8'd190;  #10 
a = 8'd196; b = 8'd191;  #10 
a = 8'd196; b = 8'd192;  #10 
a = 8'd196; b = 8'd193;  #10 
a = 8'd196; b = 8'd194;  #10 
a = 8'd196; b = 8'd195;  #10 
a = 8'd196; b = 8'd196;  #10 
a = 8'd196; b = 8'd197;  #10 
a = 8'd196; b = 8'd198;  #10 
a = 8'd196; b = 8'd199;  #10 
a = 8'd196; b = 8'd200;  #10 
a = 8'd196; b = 8'd201;  #10 
a = 8'd196; b = 8'd202;  #10 
a = 8'd196; b = 8'd203;  #10 
a = 8'd196; b = 8'd204;  #10 
a = 8'd196; b = 8'd205;  #10 
a = 8'd196; b = 8'd206;  #10 
a = 8'd196; b = 8'd207;  #10 
a = 8'd196; b = 8'd208;  #10 
a = 8'd196; b = 8'd209;  #10 
a = 8'd196; b = 8'd210;  #10 
a = 8'd196; b = 8'd211;  #10 
a = 8'd196; b = 8'd212;  #10 
a = 8'd196; b = 8'd213;  #10 
a = 8'd196; b = 8'd214;  #10 
a = 8'd196; b = 8'd215;  #10 
a = 8'd196; b = 8'd216;  #10 
a = 8'd196; b = 8'd217;  #10 
a = 8'd196; b = 8'd218;  #10 
a = 8'd196; b = 8'd219;  #10 
a = 8'd196; b = 8'd220;  #10 
a = 8'd196; b = 8'd221;  #10 
a = 8'd196; b = 8'd222;  #10 
a = 8'd196; b = 8'd223;  #10 
a = 8'd196; b = 8'd224;  #10 
a = 8'd196; b = 8'd225;  #10 
a = 8'd196; b = 8'd226;  #10 
a = 8'd196; b = 8'd227;  #10 
a = 8'd196; b = 8'd228;  #10 
a = 8'd196; b = 8'd229;  #10 
a = 8'd196; b = 8'd230;  #10 
a = 8'd196; b = 8'd231;  #10 
a = 8'd196; b = 8'd232;  #10 
a = 8'd196; b = 8'd233;  #10 
a = 8'd196; b = 8'd234;  #10 
a = 8'd196; b = 8'd235;  #10 
a = 8'd196; b = 8'd236;  #10 
a = 8'd196; b = 8'd237;  #10 
a = 8'd196; b = 8'd238;  #10 
a = 8'd196; b = 8'd239;  #10 
a = 8'd196; b = 8'd240;  #10 
a = 8'd196; b = 8'd241;  #10 
a = 8'd196; b = 8'd242;  #10 
a = 8'd196; b = 8'd243;  #10 
a = 8'd196; b = 8'd244;  #10 
a = 8'd196; b = 8'd245;  #10 
a = 8'd196; b = 8'd246;  #10 
a = 8'd196; b = 8'd247;  #10 
a = 8'd196; b = 8'd248;  #10 
a = 8'd196; b = 8'd249;  #10 
a = 8'd196; b = 8'd250;  #10 
a = 8'd196; b = 8'd251;  #10 
a = 8'd196; b = 8'd252;  #10 
a = 8'd196; b = 8'd253;  #10 
a = 8'd196; b = 8'd254;  #10 
a = 8'd196; b = 8'd255;  #10 
a = 8'd197; b = 8'd0;  #10 
a = 8'd197; b = 8'd1;  #10 
a = 8'd197; b = 8'd2;  #10 
a = 8'd197; b = 8'd3;  #10 
a = 8'd197; b = 8'd4;  #10 
a = 8'd197; b = 8'd5;  #10 
a = 8'd197; b = 8'd6;  #10 
a = 8'd197; b = 8'd7;  #10 
a = 8'd197; b = 8'd8;  #10 
a = 8'd197; b = 8'd9;  #10 
a = 8'd197; b = 8'd10;  #10 
a = 8'd197; b = 8'd11;  #10 
a = 8'd197; b = 8'd12;  #10 
a = 8'd197; b = 8'd13;  #10 
a = 8'd197; b = 8'd14;  #10 
a = 8'd197; b = 8'd15;  #10 
a = 8'd197; b = 8'd16;  #10 
a = 8'd197; b = 8'd17;  #10 
a = 8'd197; b = 8'd18;  #10 
a = 8'd197; b = 8'd19;  #10 
a = 8'd197; b = 8'd20;  #10 
a = 8'd197; b = 8'd21;  #10 
a = 8'd197; b = 8'd22;  #10 
a = 8'd197; b = 8'd23;  #10 
a = 8'd197; b = 8'd24;  #10 
a = 8'd197; b = 8'd25;  #10 
a = 8'd197; b = 8'd26;  #10 
a = 8'd197; b = 8'd27;  #10 
a = 8'd197; b = 8'd28;  #10 
a = 8'd197; b = 8'd29;  #10 
a = 8'd197; b = 8'd30;  #10 
a = 8'd197; b = 8'd31;  #10 
a = 8'd197; b = 8'd32;  #10 
a = 8'd197; b = 8'd33;  #10 
a = 8'd197; b = 8'd34;  #10 
a = 8'd197; b = 8'd35;  #10 
a = 8'd197; b = 8'd36;  #10 
a = 8'd197; b = 8'd37;  #10 
a = 8'd197; b = 8'd38;  #10 
a = 8'd197; b = 8'd39;  #10 
a = 8'd197; b = 8'd40;  #10 
a = 8'd197; b = 8'd41;  #10 
a = 8'd197; b = 8'd42;  #10 
a = 8'd197; b = 8'd43;  #10 
a = 8'd197; b = 8'd44;  #10 
a = 8'd197; b = 8'd45;  #10 
a = 8'd197; b = 8'd46;  #10 
a = 8'd197; b = 8'd47;  #10 
a = 8'd197; b = 8'd48;  #10 
a = 8'd197; b = 8'd49;  #10 
a = 8'd197; b = 8'd50;  #10 
a = 8'd197; b = 8'd51;  #10 
a = 8'd197; b = 8'd52;  #10 
a = 8'd197; b = 8'd53;  #10 
a = 8'd197; b = 8'd54;  #10 
a = 8'd197; b = 8'd55;  #10 
a = 8'd197; b = 8'd56;  #10 
a = 8'd197; b = 8'd57;  #10 
a = 8'd197; b = 8'd58;  #10 
a = 8'd197; b = 8'd59;  #10 
a = 8'd197; b = 8'd60;  #10 
a = 8'd197; b = 8'd61;  #10 
a = 8'd197; b = 8'd62;  #10 
a = 8'd197; b = 8'd63;  #10 
a = 8'd197; b = 8'd64;  #10 
a = 8'd197; b = 8'd65;  #10 
a = 8'd197; b = 8'd66;  #10 
a = 8'd197; b = 8'd67;  #10 
a = 8'd197; b = 8'd68;  #10 
a = 8'd197; b = 8'd69;  #10 
a = 8'd197; b = 8'd70;  #10 
a = 8'd197; b = 8'd71;  #10 
a = 8'd197; b = 8'd72;  #10 
a = 8'd197; b = 8'd73;  #10 
a = 8'd197; b = 8'd74;  #10 
a = 8'd197; b = 8'd75;  #10 
a = 8'd197; b = 8'd76;  #10 
a = 8'd197; b = 8'd77;  #10 
a = 8'd197; b = 8'd78;  #10 
a = 8'd197; b = 8'd79;  #10 
a = 8'd197; b = 8'd80;  #10 
a = 8'd197; b = 8'd81;  #10 
a = 8'd197; b = 8'd82;  #10 
a = 8'd197; b = 8'd83;  #10 
a = 8'd197; b = 8'd84;  #10 
a = 8'd197; b = 8'd85;  #10 
a = 8'd197; b = 8'd86;  #10 
a = 8'd197; b = 8'd87;  #10 
a = 8'd197; b = 8'd88;  #10 
a = 8'd197; b = 8'd89;  #10 
a = 8'd197; b = 8'd90;  #10 
a = 8'd197; b = 8'd91;  #10 
a = 8'd197; b = 8'd92;  #10 
a = 8'd197; b = 8'd93;  #10 
a = 8'd197; b = 8'd94;  #10 
a = 8'd197; b = 8'd95;  #10 
a = 8'd197; b = 8'd96;  #10 
a = 8'd197; b = 8'd97;  #10 
a = 8'd197; b = 8'd98;  #10 
a = 8'd197; b = 8'd99;  #10 
a = 8'd197; b = 8'd100;  #10 
a = 8'd197; b = 8'd101;  #10 
a = 8'd197; b = 8'd102;  #10 
a = 8'd197; b = 8'd103;  #10 
a = 8'd197; b = 8'd104;  #10 
a = 8'd197; b = 8'd105;  #10 
a = 8'd197; b = 8'd106;  #10 
a = 8'd197; b = 8'd107;  #10 
a = 8'd197; b = 8'd108;  #10 
a = 8'd197; b = 8'd109;  #10 
a = 8'd197; b = 8'd110;  #10 
a = 8'd197; b = 8'd111;  #10 
a = 8'd197; b = 8'd112;  #10 
a = 8'd197; b = 8'd113;  #10 
a = 8'd197; b = 8'd114;  #10 
a = 8'd197; b = 8'd115;  #10 
a = 8'd197; b = 8'd116;  #10 
a = 8'd197; b = 8'd117;  #10 
a = 8'd197; b = 8'd118;  #10 
a = 8'd197; b = 8'd119;  #10 
a = 8'd197; b = 8'd120;  #10 
a = 8'd197; b = 8'd121;  #10 
a = 8'd197; b = 8'd122;  #10 
a = 8'd197; b = 8'd123;  #10 
a = 8'd197; b = 8'd124;  #10 
a = 8'd197; b = 8'd125;  #10 
a = 8'd197; b = 8'd126;  #10 
a = 8'd197; b = 8'd127;  #10 
a = 8'd197; b = 8'd128;  #10 
a = 8'd197; b = 8'd129;  #10 
a = 8'd197; b = 8'd130;  #10 
a = 8'd197; b = 8'd131;  #10 
a = 8'd197; b = 8'd132;  #10 
a = 8'd197; b = 8'd133;  #10 
a = 8'd197; b = 8'd134;  #10 
a = 8'd197; b = 8'd135;  #10 
a = 8'd197; b = 8'd136;  #10 
a = 8'd197; b = 8'd137;  #10 
a = 8'd197; b = 8'd138;  #10 
a = 8'd197; b = 8'd139;  #10 
a = 8'd197; b = 8'd140;  #10 
a = 8'd197; b = 8'd141;  #10 
a = 8'd197; b = 8'd142;  #10 
a = 8'd197; b = 8'd143;  #10 
a = 8'd197; b = 8'd144;  #10 
a = 8'd197; b = 8'd145;  #10 
a = 8'd197; b = 8'd146;  #10 
a = 8'd197; b = 8'd147;  #10 
a = 8'd197; b = 8'd148;  #10 
a = 8'd197; b = 8'd149;  #10 
a = 8'd197; b = 8'd150;  #10 
a = 8'd197; b = 8'd151;  #10 
a = 8'd197; b = 8'd152;  #10 
a = 8'd197; b = 8'd153;  #10 
a = 8'd197; b = 8'd154;  #10 
a = 8'd197; b = 8'd155;  #10 
a = 8'd197; b = 8'd156;  #10 
a = 8'd197; b = 8'd157;  #10 
a = 8'd197; b = 8'd158;  #10 
a = 8'd197; b = 8'd159;  #10 
a = 8'd197; b = 8'd160;  #10 
a = 8'd197; b = 8'd161;  #10 
a = 8'd197; b = 8'd162;  #10 
a = 8'd197; b = 8'd163;  #10 
a = 8'd197; b = 8'd164;  #10 
a = 8'd197; b = 8'd165;  #10 
a = 8'd197; b = 8'd166;  #10 
a = 8'd197; b = 8'd167;  #10 
a = 8'd197; b = 8'd168;  #10 
a = 8'd197; b = 8'd169;  #10 
a = 8'd197; b = 8'd170;  #10 
a = 8'd197; b = 8'd171;  #10 
a = 8'd197; b = 8'd172;  #10 
a = 8'd197; b = 8'd173;  #10 
a = 8'd197; b = 8'd174;  #10 
a = 8'd197; b = 8'd175;  #10 
a = 8'd197; b = 8'd176;  #10 
a = 8'd197; b = 8'd177;  #10 
a = 8'd197; b = 8'd178;  #10 
a = 8'd197; b = 8'd179;  #10 
a = 8'd197; b = 8'd180;  #10 
a = 8'd197; b = 8'd181;  #10 
a = 8'd197; b = 8'd182;  #10 
a = 8'd197; b = 8'd183;  #10 
a = 8'd197; b = 8'd184;  #10 
a = 8'd197; b = 8'd185;  #10 
a = 8'd197; b = 8'd186;  #10 
a = 8'd197; b = 8'd187;  #10 
a = 8'd197; b = 8'd188;  #10 
a = 8'd197; b = 8'd189;  #10 
a = 8'd197; b = 8'd190;  #10 
a = 8'd197; b = 8'd191;  #10 
a = 8'd197; b = 8'd192;  #10 
a = 8'd197; b = 8'd193;  #10 
a = 8'd197; b = 8'd194;  #10 
a = 8'd197; b = 8'd195;  #10 
a = 8'd197; b = 8'd196;  #10 
a = 8'd197; b = 8'd197;  #10 
a = 8'd197; b = 8'd198;  #10 
a = 8'd197; b = 8'd199;  #10 
a = 8'd197; b = 8'd200;  #10 
a = 8'd197; b = 8'd201;  #10 
a = 8'd197; b = 8'd202;  #10 
a = 8'd197; b = 8'd203;  #10 
a = 8'd197; b = 8'd204;  #10 
a = 8'd197; b = 8'd205;  #10 
a = 8'd197; b = 8'd206;  #10 
a = 8'd197; b = 8'd207;  #10 
a = 8'd197; b = 8'd208;  #10 
a = 8'd197; b = 8'd209;  #10 
a = 8'd197; b = 8'd210;  #10 
a = 8'd197; b = 8'd211;  #10 
a = 8'd197; b = 8'd212;  #10 
a = 8'd197; b = 8'd213;  #10 
a = 8'd197; b = 8'd214;  #10 
a = 8'd197; b = 8'd215;  #10 
a = 8'd197; b = 8'd216;  #10 
a = 8'd197; b = 8'd217;  #10 
a = 8'd197; b = 8'd218;  #10 
a = 8'd197; b = 8'd219;  #10 
a = 8'd197; b = 8'd220;  #10 
a = 8'd197; b = 8'd221;  #10 
a = 8'd197; b = 8'd222;  #10 
a = 8'd197; b = 8'd223;  #10 
a = 8'd197; b = 8'd224;  #10 
a = 8'd197; b = 8'd225;  #10 
a = 8'd197; b = 8'd226;  #10 
a = 8'd197; b = 8'd227;  #10 
a = 8'd197; b = 8'd228;  #10 
a = 8'd197; b = 8'd229;  #10 
a = 8'd197; b = 8'd230;  #10 
a = 8'd197; b = 8'd231;  #10 
a = 8'd197; b = 8'd232;  #10 
a = 8'd197; b = 8'd233;  #10 
a = 8'd197; b = 8'd234;  #10 
a = 8'd197; b = 8'd235;  #10 
a = 8'd197; b = 8'd236;  #10 
a = 8'd197; b = 8'd237;  #10 
a = 8'd197; b = 8'd238;  #10 
a = 8'd197; b = 8'd239;  #10 
a = 8'd197; b = 8'd240;  #10 
a = 8'd197; b = 8'd241;  #10 
a = 8'd197; b = 8'd242;  #10 
a = 8'd197; b = 8'd243;  #10 
a = 8'd197; b = 8'd244;  #10 
a = 8'd197; b = 8'd245;  #10 
a = 8'd197; b = 8'd246;  #10 
a = 8'd197; b = 8'd247;  #10 
a = 8'd197; b = 8'd248;  #10 
a = 8'd197; b = 8'd249;  #10 
a = 8'd197; b = 8'd250;  #10 
a = 8'd197; b = 8'd251;  #10 
a = 8'd197; b = 8'd252;  #10 
a = 8'd197; b = 8'd253;  #10 
a = 8'd197; b = 8'd254;  #10 
a = 8'd197; b = 8'd255;  #10 
a = 8'd198; b = 8'd0;  #10 
a = 8'd198; b = 8'd1;  #10 
a = 8'd198; b = 8'd2;  #10 
a = 8'd198; b = 8'd3;  #10 
a = 8'd198; b = 8'd4;  #10 
a = 8'd198; b = 8'd5;  #10 
a = 8'd198; b = 8'd6;  #10 
a = 8'd198; b = 8'd7;  #10 
a = 8'd198; b = 8'd8;  #10 
a = 8'd198; b = 8'd9;  #10 
a = 8'd198; b = 8'd10;  #10 
a = 8'd198; b = 8'd11;  #10 
a = 8'd198; b = 8'd12;  #10 
a = 8'd198; b = 8'd13;  #10 
a = 8'd198; b = 8'd14;  #10 
a = 8'd198; b = 8'd15;  #10 
a = 8'd198; b = 8'd16;  #10 
a = 8'd198; b = 8'd17;  #10 
a = 8'd198; b = 8'd18;  #10 
a = 8'd198; b = 8'd19;  #10 
a = 8'd198; b = 8'd20;  #10 
a = 8'd198; b = 8'd21;  #10 
a = 8'd198; b = 8'd22;  #10 
a = 8'd198; b = 8'd23;  #10 
a = 8'd198; b = 8'd24;  #10 
a = 8'd198; b = 8'd25;  #10 
a = 8'd198; b = 8'd26;  #10 
a = 8'd198; b = 8'd27;  #10 
a = 8'd198; b = 8'd28;  #10 
a = 8'd198; b = 8'd29;  #10 
a = 8'd198; b = 8'd30;  #10 
a = 8'd198; b = 8'd31;  #10 
a = 8'd198; b = 8'd32;  #10 
a = 8'd198; b = 8'd33;  #10 
a = 8'd198; b = 8'd34;  #10 
a = 8'd198; b = 8'd35;  #10 
a = 8'd198; b = 8'd36;  #10 
a = 8'd198; b = 8'd37;  #10 
a = 8'd198; b = 8'd38;  #10 
a = 8'd198; b = 8'd39;  #10 
a = 8'd198; b = 8'd40;  #10 
a = 8'd198; b = 8'd41;  #10 
a = 8'd198; b = 8'd42;  #10 
a = 8'd198; b = 8'd43;  #10 
a = 8'd198; b = 8'd44;  #10 
a = 8'd198; b = 8'd45;  #10 
a = 8'd198; b = 8'd46;  #10 
a = 8'd198; b = 8'd47;  #10 
a = 8'd198; b = 8'd48;  #10 
a = 8'd198; b = 8'd49;  #10 
a = 8'd198; b = 8'd50;  #10 
a = 8'd198; b = 8'd51;  #10 
a = 8'd198; b = 8'd52;  #10 
a = 8'd198; b = 8'd53;  #10 
a = 8'd198; b = 8'd54;  #10 
a = 8'd198; b = 8'd55;  #10 
a = 8'd198; b = 8'd56;  #10 
a = 8'd198; b = 8'd57;  #10 
a = 8'd198; b = 8'd58;  #10 
a = 8'd198; b = 8'd59;  #10 
a = 8'd198; b = 8'd60;  #10 
a = 8'd198; b = 8'd61;  #10 
a = 8'd198; b = 8'd62;  #10 
a = 8'd198; b = 8'd63;  #10 
a = 8'd198; b = 8'd64;  #10 
a = 8'd198; b = 8'd65;  #10 
a = 8'd198; b = 8'd66;  #10 
a = 8'd198; b = 8'd67;  #10 
a = 8'd198; b = 8'd68;  #10 
a = 8'd198; b = 8'd69;  #10 
a = 8'd198; b = 8'd70;  #10 
a = 8'd198; b = 8'd71;  #10 
a = 8'd198; b = 8'd72;  #10 
a = 8'd198; b = 8'd73;  #10 
a = 8'd198; b = 8'd74;  #10 
a = 8'd198; b = 8'd75;  #10 
a = 8'd198; b = 8'd76;  #10 
a = 8'd198; b = 8'd77;  #10 
a = 8'd198; b = 8'd78;  #10 
a = 8'd198; b = 8'd79;  #10 
a = 8'd198; b = 8'd80;  #10 
a = 8'd198; b = 8'd81;  #10 
a = 8'd198; b = 8'd82;  #10 
a = 8'd198; b = 8'd83;  #10 
a = 8'd198; b = 8'd84;  #10 
a = 8'd198; b = 8'd85;  #10 
a = 8'd198; b = 8'd86;  #10 
a = 8'd198; b = 8'd87;  #10 
a = 8'd198; b = 8'd88;  #10 
a = 8'd198; b = 8'd89;  #10 
a = 8'd198; b = 8'd90;  #10 
a = 8'd198; b = 8'd91;  #10 
a = 8'd198; b = 8'd92;  #10 
a = 8'd198; b = 8'd93;  #10 
a = 8'd198; b = 8'd94;  #10 
a = 8'd198; b = 8'd95;  #10 
a = 8'd198; b = 8'd96;  #10 
a = 8'd198; b = 8'd97;  #10 
a = 8'd198; b = 8'd98;  #10 
a = 8'd198; b = 8'd99;  #10 
a = 8'd198; b = 8'd100;  #10 
a = 8'd198; b = 8'd101;  #10 
a = 8'd198; b = 8'd102;  #10 
a = 8'd198; b = 8'd103;  #10 
a = 8'd198; b = 8'd104;  #10 
a = 8'd198; b = 8'd105;  #10 
a = 8'd198; b = 8'd106;  #10 
a = 8'd198; b = 8'd107;  #10 
a = 8'd198; b = 8'd108;  #10 
a = 8'd198; b = 8'd109;  #10 
a = 8'd198; b = 8'd110;  #10 
a = 8'd198; b = 8'd111;  #10 
a = 8'd198; b = 8'd112;  #10 
a = 8'd198; b = 8'd113;  #10 
a = 8'd198; b = 8'd114;  #10 
a = 8'd198; b = 8'd115;  #10 
a = 8'd198; b = 8'd116;  #10 
a = 8'd198; b = 8'd117;  #10 
a = 8'd198; b = 8'd118;  #10 
a = 8'd198; b = 8'd119;  #10 
a = 8'd198; b = 8'd120;  #10 
a = 8'd198; b = 8'd121;  #10 
a = 8'd198; b = 8'd122;  #10 
a = 8'd198; b = 8'd123;  #10 
a = 8'd198; b = 8'd124;  #10 
a = 8'd198; b = 8'd125;  #10 
a = 8'd198; b = 8'd126;  #10 
a = 8'd198; b = 8'd127;  #10 
a = 8'd198; b = 8'd128;  #10 
a = 8'd198; b = 8'd129;  #10 
a = 8'd198; b = 8'd130;  #10 
a = 8'd198; b = 8'd131;  #10 
a = 8'd198; b = 8'd132;  #10 
a = 8'd198; b = 8'd133;  #10 
a = 8'd198; b = 8'd134;  #10 
a = 8'd198; b = 8'd135;  #10 
a = 8'd198; b = 8'd136;  #10 
a = 8'd198; b = 8'd137;  #10 
a = 8'd198; b = 8'd138;  #10 
a = 8'd198; b = 8'd139;  #10 
a = 8'd198; b = 8'd140;  #10 
a = 8'd198; b = 8'd141;  #10 
a = 8'd198; b = 8'd142;  #10 
a = 8'd198; b = 8'd143;  #10 
a = 8'd198; b = 8'd144;  #10 
a = 8'd198; b = 8'd145;  #10 
a = 8'd198; b = 8'd146;  #10 
a = 8'd198; b = 8'd147;  #10 
a = 8'd198; b = 8'd148;  #10 
a = 8'd198; b = 8'd149;  #10 
a = 8'd198; b = 8'd150;  #10 
a = 8'd198; b = 8'd151;  #10 
a = 8'd198; b = 8'd152;  #10 
a = 8'd198; b = 8'd153;  #10 
a = 8'd198; b = 8'd154;  #10 
a = 8'd198; b = 8'd155;  #10 
a = 8'd198; b = 8'd156;  #10 
a = 8'd198; b = 8'd157;  #10 
a = 8'd198; b = 8'd158;  #10 
a = 8'd198; b = 8'd159;  #10 
a = 8'd198; b = 8'd160;  #10 
a = 8'd198; b = 8'd161;  #10 
a = 8'd198; b = 8'd162;  #10 
a = 8'd198; b = 8'd163;  #10 
a = 8'd198; b = 8'd164;  #10 
a = 8'd198; b = 8'd165;  #10 
a = 8'd198; b = 8'd166;  #10 
a = 8'd198; b = 8'd167;  #10 
a = 8'd198; b = 8'd168;  #10 
a = 8'd198; b = 8'd169;  #10 
a = 8'd198; b = 8'd170;  #10 
a = 8'd198; b = 8'd171;  #10 
a = 8'd198; b = 8'd172;  #10 
a = 8'd198; b = 8'd173;  #10 
a = 8'd198; b = 8'd174;  #10 
a = 8'd198; b = 8'd175;  #10 
a = 8'd198; b = 8'd176;  #10 
a = 8'd198; b = 8'd177;  #10 
a = 8'd198; b = 8'd178;  #10 
a = 8'd198; b = 8'd179;  #10 
a = 8'd198; b = 8'd180;  #10 
a = 8'd198; b = 8'd181;  #10 
a = 8'd198; b = 8'd182;  #10 
a = 8'd198; b = 8'd183;  #10 
a = 8'd198; b = 8'd184;  #10 
a = 8'd198; b = 8'd185;  #10 
a = 8'd198; b = 8'd186;  #10 
a = 8'd198; b = 8'd187;  #10 
a = 8'd198; b = 8'd188;  #10 
a = 8'd198; b = 8'd189;  #10 
a = 8'd198; b = 8'd190;  #10 
a = 8'd198; b = 8'd191;  #10 
a = 8'd198; b = 8'd192;  #10 
a = 8'd198; b = 8'd193;  #10 
a = 8'd198; b = 8'd194;  #10 
a = 8'd198; b = 8'd195;  #10 
a = 8'd198; b = 8'd196;  #10 
a = 8'd198; b = 8'd197;  #10 
a = 8'd198; b = 8'd198;  #10 
a = 8'd198; b = 8'd199;  #10 
a = 8'd198; b = 8'd200;  #10 
a = 8'd198; b = 8'd201;  #10 
a = 8'd198; b = 8'd202;  #10 
a = 8'd198; b = 8'd203;  #10 
a = 8'd198; b = 8'd204;  #10 
a = 8'd198; b = 8'd205;  #10 
a = 8'd198; b = 8'd206;  #10 
a = 8'd198; b = 8'd207;  #10 
a = 8'd198; b = 8'd208;  #10 
a = 8'd198; b = 8'd209;  #10 
a = 8'd198; b = 8'd210;  #10 
a = 8'd198; b = 8'd211;  #10 
a = 8'd198; b = 8'd212;  #10 
a = 8'd198; b = 8'd213;  #10 
a = 8'd198; b = 8'd214;  #10 
a = 8'd198; b = 8'd215;  #10 
a = 8'd198; b = 8'd216;  #10 
a = 8'd198; b = 8'd217;  #10 
a = 8'd198; b = 8'd218;  #10 
a = 8'd198; b = 8'd219;  #10 
a = 8'd198; b = 8'd220;  #10 
a = 8'd198; b = 8'd221;  #10 
a = 8'd198; b = 8'd222;  #10 
a = 8'd198; b = 8'd223;  #10 
a = 8'd198; b = 8'd224;  #10 
a = 8'd198; b = 8'd225;  #10 
a = 8'd198; b = 8'd226;  #10 
a = 8'd198; b = 8'd227;  #10 
a = 8'd198; b = 8'd228;  #10 
a = 8'd198; b = 8'd229;  #10 
a = 8'd198; b = 8'd230;  #10 
a = 8'd198; b = 8'd231;  #10 
a = 8'd198; b = 8'd232;  #10 
a = 8'd198; b = 8'd233;  #10 
a = 8'd198; b = 8'd234;  #10 
a = 8'd198; b = 8'd235;  #10 
a = 8'd198; b = 8'd236;  #10 
a = 8'd198; b = 8'd237;  #10 
a = 8'd198; b = 8'd238;  #10 
a = 8'd198; b = 8'd239;  #10 
a = 8'd198; b = 8'd240;  #10 
a = 8'd198; b = 8'd241;  #10 
a = 8'd198; b = 8'd242;  #10 
a = 8'd198; b = 8'd243;  #10 
a = 8'd198; b = 8'd244;  #10 
a = 8'd198; b = 8'd245;  #10 
a = 8'd198; b = 8'd246;  #10 
a = 8'd198; b = 8'd247;  #10 
a = 8'd198; b = 8'd248;  #10 
a = 8'd198; b = 8'd249;  #10 
a = 8'd198; b = 8'd250;  #10 
a = 8'd198; b = 8'd251;  #10 
a = 8'd198; b = 8'd252;  #10 
a = 8'd198; b = 8'd253;  #10 
a = 8'd198; b = 8'd254;  #10 
a = 8'd198; b = 8'd255;  #10 
a = 8'd199; b = 8'd0;  #10 
a = 8'd199; b = 8'd1;  #10 
a = 8'd199; b = 8'd2;  #10 
a = 8'd199; b = 8'd3;  #10 
a = 8'd199; b = 8'd4;  #10 
a = 8'd199; b = 8'd5;  #10 
a = 8'd199; b = 8'd6;  #10 
a = 8'd199; b = 8'd7;  #10 
a = 8'd199; b = 8'd8;  #10 
a = 8'd199; b = 8'd9;  #10 
a = 8'd199; b = 8'd10;  #10 
a = 8'd199; b = 8'd11;  #10 
a = 8'd199; b = 8'd12;  #10 
a = 8'd199; b = 8'd13;  #10 
a = 8'd199; b = 8'd14;  #10 
a = 8'd199; b = 8'd15;  #10 
a = 8'd199; b = 8'd16;  #10 
a = 8'd199; b = 8'd17;  #10 
a = 8'd199; b = 8'd18;  #10 
a = 8'd199; b = 8'd19;  #10 
a = 8'd199; b = 8'd20;  #10 
a = 8'd199; b = 8'd21;  #10 
a = 8'd199; b = 8'd22;  #10 
a = 8'd199; b = 8'd23;  #10 
a = 8'd199; b = 8'd24;  #10 
a = 8'd199; b = 8'd25;  #10 
a = 8'd199; b = 8'd26;  #10 
a = 8'd199; b = 8'd27;  #10 
a = 8'd199; b = 8'd28;  #10 
a = 8'd199; b = 8'd29;  #10 
a = 8'd199; b = 8'd30;  #10 
a = 8'd199; b = 8'd31;  #10 
a = 8'd199; b = 8'd32;  #10 
a = 8'd199; b = 8'd33;  #10 
a = 8'd199; b = 8'd34;  #10 
a = 8'd199; b = 8'd35;  #10 
a = 8'd199; b = 8'd36;  #10 
a = 8'd199; b = 8'd37;  #10 
a = 8'd199; b = 8'd38;  #10 
a = 8'd199; b = 8'd39;  #10 
a = 8'd199; b = 8'd40;  #10 
a = 8'd199; b = 8'd41;  #10 
a = 8'd199; b = 8'd42;  #10 
a = 8'd199; b = 8'd43;  #10 
a = 8'd199; b = 8'd44;  #10 
a = 8'd199; b = 8'd45;  #10 
a = 8'd199; b = 8'd46;  #10 
a = 8'd199; b = 8'd47;  #10 
a = 8'd199; b = 8'd48;  #10 
a = 8'd199; b = 8'd49;  #10 
a = 8'd199; b = 8'd50;  #10 
a = 8'd199; b = 8'd51;  #10 
a = 8'd199; b = 8'd52;  #10 
a = 8'd199; b = 8'd53;  #10 
a = 8'd199; b = 8'd54;  #10 
a = 8'd199; b = 8'd55;  #10 
a = 8'd199; b = 8'd56;  #10 
a = 8'd199; b = 8'd57;  #10 
a = 8'd199; b = 8'd58;  #10 
a = 8'd199; b = 8'd59;  #10 
a = 8'd199; b = 8'd60;  #10 
a = 8'd199; b = 8'd61;  #10 
a = 8'd199; b = 8'd62;  #10 
a = 8'd199; b = 8'd63;  #10 
a = 8'd199; b = 8'd64;  #10 
a = 8'd199; b = 8'd65;  #10 
a = 8'd199; b = 8'd66;  #10 
a = 8'd199; b = 8'd67;  #10 
a = 8'd199; b = 8'd68;  #10 
a = 8'd199; b = 8'd69;  #10 
a = 8'd199; b = 8'd70;  #10 
a = 8'd199; b = 8'd71;  #10 
a = 8'd199; b = 8'd72;  #10 
a = 8'd199; b = 8'd73;  #10 
a = 8'd199; b = 8'd74;  #10 
a = 8'd199; b = 8'd75;  #10 
a = 8'd199; b = 8'd76;  #10 
a = 8'd199; b = 8'd77;  #10 
a = 8'd199; b = 8'd78;  #10 
a = 8'd199; b = 8'd79;  #10 
a = 8'd199; b = 8'd80;  #10 
a = 8'd199; b = 8'd81;  #10 
a = 8'd199; b = 8'd82;  #10 
a = 8'd199; b = 8'd83;  #10 
a = 8'd199; b = 8'd84;  #10 
a = 8'd199; b = 8'd85;  #10 
a = 8'd199; b = 8'd86;  #10 
a = 8'd199; b = 8'd87;  #10 
a = 8'd199; b = 8'd88;  #10 
a = 8'd199; b = 8'd89;  #10 
a = 8'd199; b = 8'd90;  #10 
a = 8'd199; b = 8'd91;  #10 
a = 8'd199; b = 8'd92;  #10 
a = 8'd199; b = 8'd93;  #10 
a = 8'd199; b = 8'd94;  #10 
a = 8'd199; b = 8'd95;  #10 
a = 8'd199; b = 8'd96;  #10 
a = 8'd199; b = 8'd97;  #10 
a = 8'd199; b = 8'd98;  #10 
a = 8'd199; b = 8'd99;  #10 
a = 8'd199; b = 8'd100;  #10 
a = 8'd199; b = 8'd101;  #10 
a = 8'd199; b = 8'd102;  #10 
a = 8'd199; b = 8'd103;  #10 
a = 8'd199; b = 8'd104;  #10 
a = 8'd199; b = 8'd105;  #10 
a = 8'd199; b = 8'd106;  #10 
a = 8'd199; b = 8'd107;  #10 
a = 8'd199; b = 8'd108;  #10 
a = 8'd199; b = 8'd109;  #10 
a = 8'd199; b = 8'd110;  #10 
a = 8'd199; b = 8'd111;  #10 
a = 8'd199; b = 8'd112;  #10 
a = 8'd199; b = 8'd113;  #10 
a = 8'd199; b = 8'd114;  #10 
a = 8'd199; b = 8'd115;  #10 
a = 8'd199; b = 8'd116;  #10 
a = 8'd199; b = 8'd117;  #10 
a = 8'd199; b = 8'd118;  #10 
a = 8'd199; b = 8'd119;  #10 
a = 8'd199; b = 8'd120;  #10 
a = 8'd199; b = 8'd121;  #10 
a = 8'd199; b = 8'd122;  #10 
a = 8'd199; b = 8'd123;  #10 
a = 8'd199; b = 8'd124;  #10 
a = 8'd199; b = 8'd125;  #10 
a = 8'd199; b = 8'd126;  #10 
a = 8'd199; b = 8'd127;  #10 
a = 8'd199; b = 8'd128;  #10 
a = 8'd199; b = 8'd129;  #10 
a = 8'd199; b = 8'd130;  #10 
a = 8'd199; b = 8'd131;  #10 
a = 8'd199; b = 8'd132;  #10 
a = 8'd199; b = 8'd133;  #10 
a = 8'd199; b = 8'd134;  #10 
a = 8'd199; b = 8'd135;  #10 
a = 8'd199; b = 8'd136;  #10 
a = 8'd199; b = 8'd137;  #10 
a = 8'd199; b = 8'd138;  #10 
a = 8'd199; b = 8'd139;  #10 
a = 8'd199; b = 8'd140;  #10 
a = 8'd199; b = 8'd141;  #10 
a = 8'd199; b = 8'd142;  #10 
a = 8'd199; b = 8'd143;  #10 
a = 8'd199; b = 8'd144;  #10 
a = 8'd199; b = 8'd145;  #10 
a = 8'd199; b = 8'd146;  #10 
a = 8'd199; b = 8'd147;  #10 
a = 8'd199; b = 8'd148;  #10 
a = 8'd199; b = 8'd149;  #10 
a = 8'd199; b = 8'd150;  #10 
a = 8'd199; b = 8'd151;  #10 
a = 8'd199; b = 8'd152;  #10 
a = 8'd199; b = 8'd153;  #10 
a = 8'd199; b = 8'd154;  #10 
a = 8'd199; b = 8'd155;  #10 
a = 8'd199; b = 8'd156;  #10 
a = 8'd199; b = 8'd157;  #10 
a = 8'd199; b = 8'd158;  #10 
a = 8'd199; b = 8'd159;  #10 
a = 8'd199; b = 8'd160;  #10 
a = 8'd199; b = 8'd161;  #10 
a = 8'd199; b = 8'd162;  #10 
a = 8'd199; b = 8'd163;  #10 
a = 8'd199; b = 8'd164;  #10 
a = 8'd199; b = 8'd165;  #10 
a = 8'd199; b = 8'd166;  #10 
a = 8'd199; b = 8'd167;  #10 
a = 8'd199; b = 8'd168;  #10 
a = 8'd199; b = 8'd169;  #10 
a = 8'd199; b = 8'd170;  #10 
a = 8'd199; b = 8'd171;  #10 
a = 8'd199; b = 8'd172;  #10 
a = 8'd199; b = 8'd173;  #10 
a = 8'd199; b = 8'd174;  #10 
a = 8'd199; b = 8'd175;  #10 
a = 8'd199; b = 8'd176;  #10 
a = 8'd199; b = 8'd177;  #10 
a = 8'd199; b = 8'd178;  #10 
a = 8'd199; b = 8'd179;  #10 
a = 8'd199; b = 8'd180;  #10 
a = 8'd199; b = 8'd181;  #10 
a = 8'd199; b = 8'd182;  #10 
a = 8'd199; b = 8'd183;  #10 
a = 8'd199; b = 8'd184;  #10 
a = 8'd199; b = 8'd185;  #10 
a = 8'd199; b = 8'd186;  #10 
a = 8'd199; b = 8'd187;  #10 
a = 8'd199; b = 8'd188;  #10 
a = 8'd199; b = 8'd189;  #10 
a = 8'd199; b = 8'd190;  #10 
a = 8'd199; b = 8'd191;  #10 
a = 8'd199; b = 8'd192;  #10 
a = 8'd199; b = 8'd193;  #10 
a = 8'd199; b = 8'd194;  #10 
a = 8'd199; b = 8'd195;  #10 
a = 8'd199; b = 8'd196;  #10 
a = 8'd199; b = 8'd197;  #10 
a = 8'd199; b = 8'd198;  #10 
a = 8'd199; b = 8'd199;  #10 
a = 8'd199; b = 8'd200;  #10 
a = 8'd199; b = 8'd201;  #10 
a = 8'd199; b = 8'd202;  #10 
a = 8'd199; b = 8'd203;  #10 
a = 8'd199; b = 8'd204;  #10 
a = 8'd199; b = 8'd205;  #10 
a = 8'd199; b = 8'd206;  #10 
a = 8'd199; b = 8'd207;  #10 
a = 8'd199; b = 8'd208;  #10 
a = 8'd199; b = 8'd209;  #10 
a = 8'd199; b = 8'd210;  #10 
a = 8'd199; b = 8'd211;  #10 
a = 8'd199; b = 8'd212;  #10 
a = 8'd199; b = 8'd213;  #10 
a = 8'd199; b = 8'd214;  #10 
a = 8'd199; b = 8'd215;  #10 
a = 8'd199; b = 8'd216;  #10 
a = 8'd199; b = 8'd217;  #10 
a = 8'd199; b = 8'd218;  #10 
a = 8'd199; b = 8'd219;  #10 
a = 8'd199; b = 8'd220;  #10 
a = 8'd199; b = 8'd221;  #10 
a = 8'd199; b = 8'd222;  #10 
a = 8'd199; b = 8'd223;  #10 
a = 8'd199; b = 8'd224;  #10 
a = 8'd199; b = 8'd225;  #10 
a = 8'd199; b = 8'd226;  #10 
a = 8'd199; b = 8'd227;  #10 
a = 8'd199; b = 8'd228;  #10 
a = 8'd199; b = 8'd229;  #10 
a = 8'd199; b = 8'd230;  #10 
a = 8'd199; b = 8'd231;  #10 
a = 8'd199; b = 8'd232;  #10 
a = 8'd199; b = 8'd233;  #10 
a = 8'd199; b = 8'd234;  #10 
a = 8'd199; b = 8'd235;  #10 
a = 8'd199; b = 8'd236;  #10 
a = 8'd199; b = 8'd237;  #10 
a = 8'd199; b = 8'd238;  #10 
a = 8'd199; b = 8'd239;  #10 
a = 8'd199; b = 8'd240;  #10 
a = 8'd199; b = 8'd241;  #10 
a = 8'd199; b = 8'd242;  #10 
a = 8'd199; b = 8'd243;  #10 
a = 8'd199; b = 8'd244;  #10 
a = 8'd199; b = 8'd245;  #10 
a = 8'd199; b = 8'd246;  #10 
a = 8'd199; b = 8'd247;  #10 
a = 8'd199; b = 8'd248;  #10 
a = 8'd199; b = 8'd249;  #10 
a = 8'd199; b = 8'd250;  #10 
a = 8'd199; b = 8'd251;  #10 
a = 8'd199; b = 8'd252;  #10 
a = 8'd199; b = 8'd253;  #10 
a = 8'd199; b = 8'd254;  #10 
a = 8'd199; b = 8'd255;  #10 
a = 8'd200; b = 8'd0;  #10 
a = 8'd200; b = 8'd1;  #10 
a = 8'd200; b = 8'd2;  #10 
a = 8'd200; b = 8'd3;  #10 
a = 8'd200; b = 8'd4;  #10 
a = 8'd200; b = 8'd5;  #10 
a = 8'd200; b = 8'd6;  #10 
a = 8'd200; b = 8'd7;  #10 
a = 8'd200; b = 8'd8;  #10 
a = 8'd200; b = 8'd9;  #10 
a = 8'd200; b = 8'd10;  #10 
a = 8'd200; b = 8'd11;  #10 
a = 8'd200; b = 8'd12;  #10 
a = 8'd200; b = 8'd13;  #10 
a = 8'd200; b = 8'd14;  #10 
a = 8'd200; b = 8'd15;  #10 
a = 8'd200; b = 8'd16;  #10 
a = 8'd200; b = 8'd17;  #10 
a = 8'd200; b = 8'd18;  #10 
a = 8'd200; b = 8'd19;  #10 
a = 8'd200; b = 8'd20;  #10 
a = 8'd200; b = 8'd21;  #10 
a = 8'd200; b = 8'd22;  #10 
a = 8'd200; b = 8'd23;  #10 
a = 8'd200; b = 8'd24;  #10 
a = 8'd200; b = 8'd25;  #10 
a = 8'd200; b = 8'd26;  #10 
a = 8'd200; b = 8'd27;  #10 
a = 8'd200; b = 8'd28;  #10 
a = 8'd200; b = 8'd29;  #10 
a = 8'd200; b = 8'd30;  #10 
a = 8'd200; b = 8'd31;  #10 
a = 8'd200; b = 8'd32;  #10 
a = 8'd200; b = 8'd33;  #10 
a = 8'd200; b = 8'd34;  #10 
a = 8'd200; b = 8'd35;  #10 
a = 8'd200; b = 8'd36;  #10 
a = 8'd200; b = 8'd37;  #10 
a = 8'd200; b = 8'd38;  #10 
a = 8'd200; b = 8'd39;  #10 
a = 8'd200; b = 8'd40;  #10 
a = 8'd200; b = 8'd41;  #10 
a = 8'd200; b = 8'd42;  #10 
a = 8'd200; b = 8'd43;  #10 
a = 8'd200; b = 8'd44;  #10 
a = 8'd200; b = 8'd45;  #10 
a = 8'd200; b = 8'd46;  #10 
a = 8'd200; b = 8'd47;  #10 
a = 8'd200; b = 8'd48;  #10 
a = 8'd200; b = 8'd49;  #10 
a = 8'd200; b = 8'd50;  #10 
a = 8'd200; b = 8'd51;  #10 
a = 8'd200; b = 8'd52;  #10 
a = 8'd200; b = 8'd53;  #10 
a = 8'd200; b = 8'd54;  #10 
a = 8'd200; b = 8'd55;  #10 
a = 8'd200; b = 8'd56;  #10 
a = 8'd200; b = 8'd57;  #10 
a = 8'd200; b = 8'd58;  #10 
a = 8'd200; b = 8'd59;  #10 
a = 8'd200; b = 8'd60;  #10 
a = 8'd200; b = 8'd61;  #10 
a = 8'd200; b = 8'd62;  #10 
a = 8'd200; b = 8'd63;  #10 
a = 8'd200; b = 8'd64;  #10 
a = 8'd200; b = 8'd65;  #10 
a = 8'd200; b = 8'd66;  #10 
a = 8'd200; b = 8'd67;  #10 
a = 8'd200; b = 8'd68;  #10 
a = 8'd200; b = 8'd69;  #10 
a = 8'd200; b = 8'd70;  #10 
a = 8'd200; b = 8'd71;  #10 
a = 8'd200; b = 8'd72;  #10 
a = 8'd200; b = 8'd73;  #10 
a = 8'd200; b = 8'd74;  #10 
a = 8'd200; b = 8'd75;  #10 
a = 8'd200; b = 8'd76;  #10 
a = 8'd200; b = 8'd77;  #10 
a = 8'd200; b = 8'd78;  #10 
a = 8'd200; b = 8'd79;  #10 
a = 8'd200; b = 8'd80;  #10 
a = 8'd200; b = 8'd81;  #10 
a = 8'd200; b = 8'd82;  #10 
a = 8'd200; b = 8'd83;  #10 
a = 8'd200; b = 8'd84;  #10 
a = 8'd200; b = 8'd85;  #10 
a = 8'd200; b = 8'd86;  #10 
a = 8'd200; b = 8'd87;  #10 
a = 8'd200; b = 8'd88;  #10 
a = 8'd200; b = 8'd89;  #10 
a = 8'd200; b = 8'd90;  #10 
a = 8'd200; b = 8'd91;  #10 
a = 8'd200; b = 8'd92;  #10 
a = 8'd200; b = 8'd93;  #10 
a = 8'd200; b = 8'd94;  #10 
a = 8'd200; b = 8'd95;  #10 
a = 8'd200; b = 8'd96;  #10 
a = 8'd200; b = 8'd97;  #10 
a = 8'd200; b = 8'd98;  #10 
a = 8'd200; b = 8'd99;  #10 
a = 8'd200; b = 8'd100;  #10 
a = 8'd200; b = 8'd101;  #10 
a = 8'd200; b = 8'd102;  #10 
a = 8'd200; b = 8'd103;  #10 
a = 8'd200; b = 8'd104;  #10 
a = 8'd200; b = 8'd105;  #10 
a = 8'd200; b = 8'd106;  #10 
a = 8'd200; b = 8'd107;  #10 
a = 8'd200; b = 8'd108;  #10 
a = 8'd200; b = 8'd109;  #10 
a = 8'd200; b = 8'd110;  #10 
a = 8'd200; b = 8'd111;  #10 
a = 8'd200; b = 8'd112;  #10 
a = 8'd200; b = 8'd113;  #10 
a = 8'd200; b = 8'd114;  #10 
a = 8'd200; b = 8'd115;  #10 
a = 8'd200; b = 8'd116;  #10 
a = 8'd200; b = 8'd117;  #10 
a = 8'd200; b = 8'd118;  #10 
a = 8'd200; b = 8'd119;  #10 
a = 8'd200; b = 8'd120;  #10 
a = 8'd200; b = 8'd121;  #10 
a = 8'd200; b = 8'd122;  #10 
a = 8'd200; b = 8'd123;  #10 
a = 8'd200; b = 8'd124;  #10 
a = 8'd200; b = 8'd125;  #10 
a = 8'd200; b = 8'd126;  #10 
a = 8'd200; b = 8'd127;  #10 
a = 8'd200; b = 8'd128;  #10 
a = 8'd200; b = 8'd129;  #10 
a = 8'd200; b = 8'd130;  #10 
a = 8'd200; b = 8'd131;  #10 
a = 8'd200; b = 8'd132;  #10 
a = 8'd200; b = 8'd133;  #10 
a = 8'd200; b = 8'd134;  #10 
a = 8'd200; b = 8'd135;  #10 
a = 8'd200; b = 8'd136;  #10 
a = 8'd200; b = 8'd137;  #10 
a = 8'd200; b = 8'd138;  #10 
a = 8'd200; b = 8'd139;  #10 
a = 8'd200; b = 8'd140;  #10 
a = 8'd200; b = 8'd141;  #10 
a = 8'd200; b = 8'd142;  #10 
a = 8'd200; b = 8'd143;  #10 
a = 8'd200; b = 8'd144;  #10 
a = 8'd200; b = 8'd145;  #10 
a = 8'd200; b = 8'd146;  #10 
a = 8'd200; b = 8'd147;  #10 
a = 8'd200; b = 8'd148;  #10 
a = 8'd200; b = 8'd149;  #10 
a = 8'd200; b = 8'd150;  #10 
a = 8'd200; b = 8'd151;  #10 
a = 8'd200; b = 8'd152;  #10 
a = 8'd200; b = 8'd153;  #10 
a = 8'd200; b = 8'd154;  #10 
a = 8'd200; b = 8'd155;  #10 
a = 8'd200; b = 8'd156;  #10 
a = 8'd200; b = 8'd157;  #10 
a = 8'd200; b = 8'd158;  #10 
a = 8'd200; b = 8'd159;  #10 
a = 8'd200; b = 8'd160;  #10 
a = 8'd200; b = 8'd161;  #10 
a = 8'd200; b = 8'd162;  #10 
a = 8'd200; b = 8'd163;  #10 
a = 8'd200; b = 8'd164;  #10 
a = 8'd200; b = 8'd165;  #10 
a = 8'd200; b = 8'd166;  #10 
a = 8'd200; b = 8'd167;  #10 
a = 8'd200; b = 8'd168;  #10 
a = 8'd200; b = 8'd169;  #10 
a = 8'd200; b = 8'd170;  #10 
a = 8'd200; b = 8'd171;  #10 
a = 8'd200; b = 8'd172;  #10 
a = 8'd200; b = 8'd173;  #10 
a = 8'd200; b = 8'd174;  #10 
a = 8'd200; b = 8'd175;  #10 
a = 8'd200; b = 8'd176;  #10 
a = 8'd200; b = 8'd177;  #10 
a = 8'd200; b = 8'd178;  #10 
a = 8'd200; b = 8'd179;  #10 
a = 8'd200; b = 8'd180;  #10 
a = 8'd200; b = 8'd181;  #10 
a = 8'd200; b = 8'd182;  #10 
a = 8'd200; b = 8'd183;  #10 
a = 8'd200; b = 8'd184;  #10 
a = 8'd200; b = 8'd185;  #10 
a = 8'd200; b = 8'd186;  #10 
a = 8'd200; b = 8'd187;  #10 
a = 8'd200; b = 8'd188;  #10 
a = 8'd200; b = 8'd189;  #10 
a = 8'd200; b = 8'd190;  #10 
a = 8'd200; b = 8'd191;  #10 
a = 8'd200; b = 8'd192;  #10 
a = 8'd200; b = 8'd193;  #10 
a = 8'd200; b = 8'd194;  #10 
a = 8'd200; b = 8'd195;  #10 
a = 8'd200; b = 8'd196;  #10 
a = 8'd200; b = 8'd197;  #10 
a = 8'd200; b = 8'd198;  #10 
a = 8'd200; b = 8'd199;  #10 
a = 8'd200; b = 8'd200;  #10 
a = 8'd200; b = 8'd201;  #10 
a = 8'd200; b = 8'd202;  #10 
a = 8'd200; b = 8'd203;  #10 
a = 8'd200; b = 8'd204;  #10 
a = 8'd200; b = 8'd205;  #10 
a = 8'd200; b = 8'd206;  #10 
a = 8'd200; b = 8'd207;  #10 
a = 8'd200; b = 8'd208;  #10 
a = 8'd200; b = 8'd209;  #10 
a = 8'd200; b = 8'd210;  #10 
a = 8'd200; b = 8'd211;  #10 
a = 8'd200; b = 8'd212;  #10 
a = 8'd200; b = 8'd213;  #10 
a = 8'd200; b = 8'd214;  #10 
a = 8'd200; b = 8'd215;  #10 
a = 8'd200; b = 8'd216;  #10 
a = 8'd200; b = 8'd217;  #10 
a = 8'd200; b = 8'd218;  #10 
a = 8'd200; b = 8'd219;  #10 
a = 8'd200; b = 8'd220;  #10 
a = 8'd200; b = 8'd221;  #10 
a = 8'd200; b = 8'd222;  #10 
a = 8'd200; b = 8'd223;  #10 
a = 8'd200; b = 8'd224;  #10 
a = 8'd200; b = 8'd225;  #10 
a = 8'd200; b = 8'd226;  #10 
a = 8'd200; b = 8'd227;  #10 
a = 8'd200; b = 8'd228;  #10 
a = 8'd200; b = 8'd229;  #10 
a = 8'd200; b = 8'd230;  #10 
a = 8'd200; b = 8'd231;  #10 
a = 8'd200; b = 8'd232;  #10 
a = 8'd200; b = 8'd233;  #10 
a = 8'd200; b = 8'd234;  #10 
a = 8'd200; b = 8'd235;  #10 
a = 8'd200; b = 8'd236;  #10 
a = 8'd200; b = 8'd237;  #10 
a = 8'd200; b = 8'd238;  #10 
a = 8'd200; b = 8'd239;  #10 
a = 8'd200; b = 8'd240;  #10 
a = 8'd200; b = 8'd241;  #10 
a = 8'd200; b = 8'd242;  #10 
a = 8'd200; b = 8'd243;  #10 
a = 8'd200; b = 8'd244;  #10 
a = 8'd200; b = 8'd245;  #10 
a = 8'd200; b = 8'd246;  #10 
a = 8'd200; b = 8'd247;  #10 
a = 8'd200; b = 8'd248;  #10 
a = 8'd200; b = 8'd249;  #10 
a = 8'd200; b = 8'd250;  #10 
a = 8'd200; b = 8'd251;  #10 
a = 8'd200; b = 8'd252;  #10 
a = 8'd200; b = 8'd253;  #10 
a = 8'd200; b = 8'd254;  #10 
a = 8'd200; b = 8'd255;  #10 
a = 8'd201; b = 8'd0;  #10 
a = 8'd201; b = 8'd1;  #10 
a = 8'd201; b = 8'd2;  #10 
a = 8'd201; b = 8'd3;  #10 
a = 8'd201; b = 8'd4;  #10 
a = 8'd201; b = 8'd5;  #10 
a = 8'd201; b = 8'd6;  #10 
a = 8'd201; b = 8'd7;  #10 
a = 8'd201; b = 8'd8;  #10 
a = 8'd201; b = 8'd9;  #10 
a = 8'd201; b = 8'd10;  #10 
a = 8'd201; b = 8'd11;  #10 
a = 8'd201; b = 8'd12;  #10 
a = 8'd201; b = 8'd13;  #10 
a = 8'd201; b = 8'd14;  #10 
a = 8'd201; b = 8'd15;  #10 
a = 8'd201; b = 8'd16;  #10 
a = 8'd201; b = 8'd17;  #10 
a = 8'd201; b = 8'd18;  #10 
a = 8'd201; b = 8'd19;  #10 
a = 8'd201; b = 8'd20;  #10 
a = 8'd201; b = 8'd21;  #10 
a = 8'd201; b = 8'd22;  #10 
a = 8'd201; b = 8'd23;  #10 
a = 8'd201; b = 8'd24;  #10 
a = 8'd201; b = 8'd25;  #10 
a = 8'd201; b = 8'd26;  #10 
a = 8'd201; b = 8'd27;  #10 
a = 8'd201; b = 8'd28;  #10 
a = 8'd201; b = 8'd29;  #10 
a = 8'd201; b = 8'd30;  #10 
a = 8'd201; b = 8'd31;  #10 
a = 8'd201; b = 8'd32;  #10 
a = 8'd201; b = 8'd33;  #10 
a = 8'd201; b = 8'd34;  #10 
a = 8'd201; b = 8'd35;  #10 
a = 8'd201; b = 8'd36;  #10 
a = 8'd201; b = 8'd37;  #10 
a = 8'd201; b = 8'd38;  #10 
a = 8'd201; b = 8'd39;  #10 
a = 8'd201; b = 8'd40;  #10 
a = 8'd201; b = 8'd41;  #10 
a = 8'd201; b = 8'd42;  #10 
a = 8'd201; b = 8'd43;  #10 
a = 8'd201; b = 8'd44;  #10 
a = 8'd201; b = 8'd45;  #10 
a = 8'd201; b = 8'd46;  #10 
a = 8'd201; b = 8'd47;  #10 
a = 8'd201; b = 8'd48;  #10 
a = 8'd201; b = 8'd49;  #10 
a = 8'd201; b = 8'd50;  #10 
a = 8'd201; b = 8'd51;  #10 
a = 8'd201; b = 8'd52;  #10 
a = 8'd201; b = 8'd53;  #10 
a = 8'd201; b = 8'd54;  #10 
a = 8'd201; b = 8'd55;  #10 
a = 8'd201; b = 8'd56;  #10 
a = 8'd201; b = 8'd57;  #10 
a = 8'd201; b = 8'd58;  #10 
a = 8'd201; b = 8'd59;  #10 
a = 8'd201; b = 8'd60;  #10 
a = 8'd201; b = 8'd61;  #10 
a = 8'd201; b = 8'd62;  #10 
a = 8'd201; b = 8'd63;  #10 
a = 8'd201; b = 8'd64;  #10 
a = 8'd201; b = 8'd65;  #10 
a = 8'd201; b = 8'd66;  #10 
a = 8'd201; b = 8'd67;  #10 
a = 8'd201; b = 8'd68;  #10 
a = 8'd201; b = 8'd69;  #10 
a = 8'd201; b = 8'd70;  #10 
a = 8'd201; b = 8'd71;  #10 
a = 8'd201; b = 8'd72;  #10 
a = 8'd201; b = 8'd73;  #10 
a = 8'd201; b = 8'd74;  #10 
a = 8'd201; b = 8'd75;  #10 
a = 8'd201; b = 8'd76;  #10 
a = 8'd201; b = 8'd77;  #10 
a = 8'd201; b = 8'd78;  #10 
a = 8'd201; b = 8'd79;  #10 
a = 8'd201; b = 8'd80;  #10 
a = 8'd201; b = 8'd81;  #10 
a = 8'd201; b = 8'd82;  #10 
a = 8'd201; b = 8'd83;  #10 
a = 8'd201; b = 8'd84;  #10 
a = 8'd201; b = 8'd85;  #10 
a = 8'd201; b = 8'd86;  #10 
a = 8'd201; b = 8'd87;  #10 
a = 8'd201; b = 8'd88;  #10 
a = 8'd201; b = 8'd89;  #10 
a = 8'd201; b = 8'd90;  #10 
a = 8'd201; b = 8'd91;  #10 
a = 8'd201; b = 8'd92;  #10 
a = 8'd201; b = 8'd93;  #10 
a = 8'd201; b = 8'd94;  #10 
a = 8'd201; b = 8'd95;  #10 
a = 8'd201; b = 8'd96;  #10 
a = 8'd201; b = 8'd97;  #10 
a = 8'd201; b = 8'd98;  #10 
a = 8'd201; b = 8'd99;  #10 
a = 8'd201; b = 8'd100;  #10 
a = 8'd201; b = 8'd101;  #10 
a = 8'd201; b = 8'd102;  #10 
a = 8'd201; b = 8'd103;  #10 
a = 8'd201; b = 8'd104;  #10 
a = 8'd201; b = 8'd105;  #10 
a = 8'd201; b = 8'd106;  #10 
a = 8'd201; b = 8'd107;  #10 
a = 8'd201; b = 8'd108;  #10 
a = 8'd201; b = 8'd109;  #10 
a = 8'd201; b = 8'd110;  #10 
a = 8'd201; b = 8'd111;  #10 
a = 8'd201; b = 8'd112;  #10 
a = 8'd201; b = 8'd113;  #10 
a = 8'd201; b = 8'd114;  #10 
a = 8'd201; b = 8'd115;  #10 
a = 8'd201; b = 8'd116;  #10 
a = 8'd201; b = 8'd117;  #10 
a = 8'd201; b = 8'd118;  #10 
a = 8'd201; b = 8'd119;  #10 
a = 8'd201; b = 8'd120;  #10 
a = 8'd201; b = 8'd121;  #10 
a = 8'd201; b = 8'd122;  #10 
a = 8'd201; b = 8'd123;  #10 
a = 8'd201; b = 8'd124;  #10 
a = 8'd201; b = 8'd125;  #10 
a = 8'd201; b = 8'd126;  #10 
a = 8'd201; b = 8'd127;  #10 
a = 8'd201; b = 8'd128;  #10 
a = 8'd201; b = 8'd129;  #10 
a = 8'd201; b = 8'd130;  #10 
a = 8'd201; b = 8'd131;  #10 
a = 8'd201; b = 8'd132;  #10 
a = 8'd201; b = 8'd133;  #10 
a = 8'd201; b = 8'd134;  #10 
a = 8'd201; b = 8'd135;  #10 
a = 8'd201; b = 8'd136;  #10 
a = 8'd201; b = 8'd137;  #10 
a = 8'd201; b = 8'd138;  #10 
a = 8'd201; b = 8'd139;  #10 
a = 8'd201; b = 8'd140;  #10 
a = 8'd201; b = 8'd141;  #10 
a = 8'd201; b = 8'd142;  #10 
a = 8'd201; b = 8'd143;  #10 
a = 8'd201; b = 8'd144;  #10 
a = 8'd201; b = 8'd145;  #10 
a = 8'd201; b = 8'd146;  #10 
a = 8'd201; b = 8'd147;  #10 
a = 8'd201; b = 8'd148;  #10 
a = 8'd201; b = 8'd149;  #10 
a = 8'd201; b = 8'd150;  #10 
a = 8'd201; b = 8'd151;  #10 
a = 8'd201; b = 8'd152;  #10 
a = 8'd201; b = 8'd153;  #10 
a = 8'd201; b = 8'd154;  #10 
a = 8'd201; b = 8'd155;  #10 
a = 8'd201; b = 8'd156;  #10 
a = 8'd201; b = 8'd157;  #10 
a = 8'd201; b = 8'd158;  #10 
a = 8'd201; b = 8'd159;  #10 
a = 8'd201; b = 8'd160;  #10 
a = 8'd201; b = 8'd161;  #10 
a = 8'd201; b = 8'd162;  #10 
a = 8'd201; b = 8'd163;  #10 
a = 8'd201; b = 8'd164;  #10 
a = 8'd201; b = 8'd165;  #10 
a = 8'd201; b = 8'd166;  #10 
a = 8'd201; b = 8'd167;  #10 
a = 8'd201; b = 8'd168;  #10 
a = 8'd201; b = 8'd169;  #10 
a = 8'd201; b = 8'd170;  #10 
a = 8'd201; b = 8'd171;  #10 
a = 8'd201; b = 8'd172;  #10 
a = 8'd201; b = 8'd173;  #10 
a = 8'd201; b = 8'd174;  #10 
a = 8'd201; b = 8'd175;  #10 
a = 8'd201; b = 8'd176;  #10 
a = 8'd201; b = 8'd177;  #10 
a = 8'd201; b = 8'd178;  #10 
a = 8'd201; b = 8'd179;  #10 
a = 8'd201; b = 8'd180;  #10 
a = 8'd201; b = 8'd181;  #10 
a = 8'd201; b = 8'd182;  #10 
a = 8'd201; b = 8'd183;  #10 
a = 8'd201; b = 8'd184;  #10 
a = 8'd201; b = 8'd185;  #10 
a = 8'd201; b = 8'd186;  #10 
a = 8'd201; b = 8'd187;  #10 
a = 8'd201; b = 8'd188;  #10 
a = 8'd201; b = 8'd189;  #10 
a = 8'd201; b = 8'd190;  #10 
a = 8'd201; b = 8'd191;  #10 
a = 8'd201; b = 8'd192;  #10 
a = 8'd201; b = 8'd193;  #10 
a = 8'd201; b = 8'd194;  #10 
a = 8'd201; b = 8'd195;  #10 
a = 8'd201; b = 8'd196;  #10 
a = 8'd201; b = 8'd197;  #10 
a = 8'd201; b = 8'd198;  #10 
a = 8'd201; b = 8'd199;  #10 
a = 8'd201; b = 8'd200;  #10 
a = 8'd201; b = 8'd201;  #10 
a = 8'd201; b = 8'd202;  #10 
a = 8'd201; b = 8'd203;  #10 
a = 8'd201; b = 8'd204;  #10 
a = 8'd201; b = 8'd205;  #10 
a = 8'd201; b = 8'd206;  #10 
a = 8'd201; b = 8'd207;  #10 
a = 8'd201; b = 8'd208;  #10 
a = 8'd201; b = 8'd209;  #10 
a = 8'd201; b = 8'd210;  #10 
a = 8'd201; b = 8'd211;  #10 
a = 8'd201; b = 8'd212;  #10 
a = 8'd201; b = 8'd213;  #10 
a = 8'd201; b = 8'd214;  #10 
a = 8'd201; b = 8'd215;  #10 
a = 8'd201; b = 8'd216;  #10 
a = 8'd201; b = 8'd217;  #10 
a = 8'd201; b = 8'd218;  #10 
a = 8'd201; b = 8'd219;  #10 
a = 8'd201; b = 8'd220;  #10 
a = 8'd201; b = 8'd221;  #10 
a = 8'd201; b = 8'd222;  #10 
a = 8'd201; b = 8'd223;  #10 
a = 8'd201; b = 8'd224;  #10 
a = 8'd201; b = 8'd225;  #10 
a = 8'd201; b = 8'd226;  #10 
a = 8'd201; b = 8'd227;  #10 
a = 8'd201; b = 8'd228;  #10 
a = 8'd201; b = 8'd229;  #10 
a = 8'd201; b = 8'd230;  #10 
a = 8'd201; b = 8'd231;  #10 
a = 8'd201; b = 8'd232;  #10 
a = 8'd201; b = 8'd233;  #10 
a = 8'd201; b = 8'd234;  #10 
a = 8'd201; b = 8'd235;  #10 
a = 8'd201; b = 8'd236;  #10 
a = 8'd201; b = 8'd237;  #10 
a = 8'd201; b = 8'd238;  #10 
a = 8'd201; b = 8'd239;  #10 
a = 8'd201; b = 8'd240;  #10 
a = 8'd201; b = 8'd241;  #10 
a = 8'd201; b = 8'd242;  #10 
a = 8'd201; b = 8'd243;  #10 
a = 8'd201; b = 8'd244;  #10 
a = 8'd201; b = 8'd245;  #10 
a = 8'd201; b = 8'd246;  #10 
a = 8'd201; b = 8'd247;  #10 
a = 8'd201; b = 8'd248;  #10 
a = 8'd201; b = 8'd249;  #10 
a = 8'd201; b = 8'd250;  #10 
a = 8'd201; b = 8'd251;  #10 
a = 8'd201; b = 8'd252;  #10 
a = 8'd201; b = 8'd253;  #10 
a = 8'd201; b = 8'd254;  #10 
a = 8'd201; b = 8'd255;  #10 
a = 8'd202; b = 8'd0;  #10 
a = 8'd202; b = 8'd1;  #10 
a = 8'd202; b = 8'd2;  #10 
a = 8'd202; b = 8'd3;  #10 
a = 8'd202; b = 8'd4;  #10 
a = 8'd202; b = 8'd5;  #10 
a = 8'd202; b = 8'd6;  #10 
a = 8'd202; b = 8'd7;  #10 
a = 8'd202; b = 8'd8;  #10 
a = 8'd202; b = 8'd9;  #10 
a = 8'd202; b = 8'd10;  #10 
a = 8'd202; b = 8'd11;  #10 
a = 8'd202; b = 8'd12;  #10 
a = 8'd202; b = 8'd13;  #10 
a = 8'd202; b = 8'd14;  #10 
a = 8'd202; b = 8'd15;  #10 
a = 8'd202; b = 8'd16;  #10 
a = 8'd202; b = 8'd17;  #10 
a = 8'd202; b = 8'd18;  #10 
a = 8'd202; b = 8'd19;  #10 
a = 8'd202; b = 8'd20;  #10 
a = 8'd202; b = 8'd21;  #10 
a = 8'd202; b = 8'd22;  #10 
a = 8'd202; b = 8'd23;  #10 
a = 8'd202; b = 8'd24;  #10 
a = 8'd202; b = 8'd25;  #10 
a = 8'd202; b = 8'd26;  #10 
a = 8'd202; b = 8'd27;  #10 
a = 8'd202; b = 8'd28;  #10 
a = 8'd202; b = 8'd29;  #10 
a = 8'd202; b = 8'd30;  #10 
a = 8'd202; b = 8'd31;  #10 
a = 8'd202; b = 8'd32;  #10 
a = 8'd202; b = 8'd33;  #10 
a = 8'd202; b = 8'd34;  #10 
a = 8'd202; b = 8'd35;  #10 
a = 8'd202; b = 8'd36;  #10 
a = 8'd202; b = 8'd37;  #10 
a = 8'd202; b = 8'd38;  #10 
a = 8'd202; b = 8'd39;  #10 
a = 8'd202; b = 8'd40;  #10 
a = 8'd202; b = 8'd41;  #10 
a = 8'd202; b = 8'd42;  #10 
a = 8'd202; b = 8'd43;  #10 
a = 8'd202; b = 8'd44;  #10 
a = 8'd202; b = 8'd45;  #10 
a = 8'd202; b = 8'd46;  #10 
a = 8'd202; b = 8'd47;  #10 
a = 8'd202; b = 8'd48;  #10 
a = 8'd202; b = 8'd49;  #10 
a = 8'd202; b = 8'd50;  #10 
a = 8'd202; b = 8'd51;  #10 
a = 8'd202; b = 8'd52;  #10 
a = 8'd202; b = 8'd53;  #10 
a = 8'd202; b = 8'd54;  #10 
a = 8'd202; b = 8'd55;  #10 
a = 8'd202; b = 8'd56;  #10 
a = 8'd202; b = 8'd57;  #10 
a = 8'd202; b = 8'd58;  #10 
a = 8'd202; b = 8'd59;  #10 
a = 8'd202; b = 8'd60;  #10 
a = 8'd202; b = 8'd61;  #10 
a = 8'd202; b = 8'd62;  #10 
a = 8'd202; b = 8'd63;  #10 
a = 8'd202; b = 8'd64;  #10 
a = 8'd202; b = 8'd65;  #10 
a = 8'd202; b = 8'd66;  #10 
a = 8'd202; b = 8'd67;  #10 
a = 8'd202; b = 8'd68;  #10 
a = 8'd202; b = 8'd69;  #10 
a = 8'd202; b = 8'd70;  #10 
a = 8'd202; b = 8'd71;  #10 
a = 8'd202; b = 8'd72;  #10 
a = 8'd202; b = 8'd73;  #10 
a = 8'd202; b = 8'd74;  #10 
a = 8'd202; b = 8'd75;  #10 
a = 8'd202; b = 8'd76;  #10 
a = 8'd202; b = 8'd77;  #10 
a = 8'd202; b = 8'd78;  #10 
a = 8'd202; b = 8'd79;  #10 
a = 8'd202; b = 8'd80;  #10 
a = 8'd202; b = 8'd81;  #10 
a = 8'd202; b = 8'd82;  #10 
a = 8'd202; b = 8'd83;  #10 
a = 8'd202; b = 8'd84;  #10 
a = 8'd202; b = 8'd85;  #10 
a = 8'd202; b = 8'd86;  #10 
a = 8'd202; b = 8'd87;  #10 
a = 8'd202; b = 8'd88;  #10 
a = 8'd202; b = 8'd89;  #10 
a = 8'd202; b = 8'd90;  #10 
a = 8'd202; b = 8'd91;  #10 
a = 8'd202; b = 8'd92;  #10 
a = 8'd202; b = 8'd93;  #10 
a = 8'd202; b = 8'd94;  #10 
a = 8'd202; b = 8'd95;  #10 
a = 8'd202; b = 8'd96;  #10 
a = 8'd202; b = 8'd97;  #10 
a = 8'd202; b = 8'd98;  #10 
a = 8'd202; b = 8'd99;  #10 
a = 8'd202; b = 8'd100;  #10 
a = 8'd202; b = 8'd101;  #10 
a = 8'd202; b = 8'd102;  #10 
a = 8'd202; b = 8'd103;  #10 
a = 8'd202; b = 8'd104;  #10 
a = 8'd202; b = 8'd105;  #10 
a = 8'd202; b = 8'd106;  #10 
a = 8'd202; b = 8'd107;  #10 
a = 8'd202; b = 8'd108;  #10 
a = 8'd202; b = 8'd109;  #10 
a = 8'd202; b = 8'd110;  #10 
a = 8'd202; b = 8'd111;  #10 
a = 8'd202; b = 8'd112;  #10 
a = 8'd202; b = 8'd113;  #10 
a = 8'd202; b = 8'd114;  #10 
a = 8'd202; b = 8'd115;  #10 
a = 8'd202; b = 8'd116;  #10 
a = 8'd202; b = 8'd117;  #10 
a = 8'd202; b = 8'd118;  #10 
a = 8'd202; b = 8'd119;  #10 
a = 8'd202; b = 8'd120;  #10 
a = 8'd202; b = 8'd121;  #10 
a = 8'd202; b = 8'd122;  #10 
a = 8'd202; b = 8'd123;  #10 
a = 8'd202; b = 8'd124;  #10 
a = 8'd202; b = 8'd125;  #10 
a = 8'd202; b = 8'd126;  #10 
a = 8'd202; b = 8'd127;  #10 
a = 8'd202; b = 8'd128;  #10 
a = 8'd202; b = 8'd129;  #10 
a = 8'd202; b = 8'd130;  #10 
a = 8'd202; b = 8'd131;  #10 
a = 8'd202; b = 8'd132;  #10 
a = 8'd202; b = 8'd133;  #10 
a = 8'd202; b = 8'd134;  #10 
a = 8'd202; b = 8'd135;  #10 
a = 8'd202; b = 8'd136;  #10 
a = 8'd202; b = 8'd137;  #10 
a = 8'd202; b = 8'd138;  #10 
a = 8'd202; b = 8'd139;  #10 
a = 8'd202; b = 8'd140;  #10 
a = 8'd202; b = 8'd141;  #10 
a = 8'd202; b = 8'd142;  #10 
a = 8'd202; b = 8'd143;  #10 
a = 8'd202; b = 8'd144;  #10 
a = 8'd202; b = 8'd145;  #10 
a = 8'd202; b = 8'd146;  #10 
a = 8'd202; b = 8'd147;  #10 
a = 8'd202; b = 8'd148;  #10 
a = 8'd202; b = 8'd149;  #10 
a = 8'd202; b = 8'd150;  #10 
a = 8'd202; b = 8'd151;  #10 
a = 8'd202; b = 8'd152;  #10 
a = 8'd202; b = 8'd153;  #10 
a = 8'd202; b = 8'd154;  #10 
a = 8'd202; b = 8'd155;  #10 
a = 8'd202; b = 8'd156;  #10 
a = 8'd202; b = 8'd157;  #10 
a = 8'd202; b = 8'd158;  #10 
a = 8'd202; b = 8'd159;  #10 
a = 8'd202; b = 8'd160;  #10 
a = 8'd202; b = 8'd161;  #10 
a = 8'd202; b = 8'd162;  #10 
a = 8'd202; b = 8'd163;  #10 
a = 8'd202; b = 8'd164;  #10 
a = 8'd202; b = 8'd165;  #10 
a = 8'd202; b = 8'd166;  #10 
a = 8'd202; b = 8'd167;  #10 
a = 8'd202; b = 8'd168;  #10 
a = 8'd202; b = 8'd169;  #10 
a = 8'd202; b = 8'd170;  #10 
a = 8'd202; b = 8'd171;  #10 
a = 8'd202; b = 8'd172;  #10 
a = 8'd202; b = 8'd173;  #10 
a = 8'd202; b = 8'd174;  #10 
a = 8'd202; b = 8'd175;  #10 
a = 8'd202; b = 8'd176;  #10 
a = 8'd202; b = 8'd177;  #10 
a = 8'd202; b = 8'd178;  #10 
a = 8'd202; b = 8'd179;  #10 
a = 8'd202; b = 8'd180;  #10 
a = 8'd202; b = 8'd181;  #10 
a = 8'd202; b = 8'd182;  #10 
a = 8'd202; b = 8'd183;  #10 
a = 8'd202; b = 8'd184;  #10 
a = 8'd202; b = 8'd185;  #10 
a = 8'd202; b = 8'd186;  #10 
a = 8'd202; b = 8'd187;  #10 
a = 8'd202; b = 8'd188;  #10 
a = 8'd202; b = 8'd189;  #10 
a = 8'd202; b = 8'd190;  #10 
a = 8'd202; b = 8'd191;  #10 
a = 8'd202; b = 8'd192;  #10 
a = 8'd202; b = 8'd193;  #10 
a = 8'd202; b = 8'd194;  #10 
a = 8'd202; b = 8'd195;  #10 
a = 8'd202; b = 8'd196;  #10 
a = 8'd202; b = 8'd197;  #10 
a = 8'd202; b = 8'd198;  #10 
a = 8'd202; b = 8'd199;  #10 
a = 8'd202; b = 8'd200;  #10 
a = 8'd202; b = 8'd201;  #10 
a = 8'd202; b = 8'd202;  #10 
a = 8'd202; b = 8'd203;  #10 
a = 8'd202; b = 8'd204;  #10 
a = 8'd202; b = 8'd205;  #10 
a = 8'd202; b = 8'd206;  #10 
a = 8'd202; b = 8'd207;  #10 
a = 8'd202; b = 8'd208;  #10 
a = 8'd202; b = 8'd209;  #10 
a = 8'd202; b = 8'd210;  #10 
a = 8'd202; b = 8'd211;  #10 
a = 8'd202; b = 8'd212;  #10 
a = 8'd202; b = 8'd213;  #10 
a = 8'd202; b = 8'd214;  #10 
a = 8'd202; b = 8'd215;  #10 
a = 8'd202; b = 8'd216;  #10 
a = 8'd202; b = 8'd217;  #10 
a = 8'd202; b = 8'd218;  #10 
a = 8'd202; b = 8'd219;  #10 
a = 8'd202; b = 8'd220;  #10 
a = 8'd202; b = 8'd221;  #10 
a = 8'd202; b = 8'd222;  #10 
a = 8'd202; b = 8'd223;  #10 
a = 8'd202; b = 8'd224;  #10 
a = 8'd202; b = 8'd225;  #10 
a = 8'd202; b = 8'd226;  #10 
a = 8'd202; b = 8'd227;  #10 
a = 8'd202; b = 8'd228;  #10 
a = 8'd202; b = 8'd229;  #10 
a = 8'd202; b = 8'd230;  #10 
a = 8'd202; b = 8'd231;  #10 
a = 8'd202; b = 8'd232;  #10 
a = 8'd202; b = 8'd233;  #10 
a = 8'd202; b = 8'd234;  #10 
a = 8'd202; b = 8'd235;  #10 
a = 8'd202; b = 8'd236;  #10 
a = 8'd202; b = 8'd237;  #10 
a = 8'd202; b = 8'd238;  #10 
a = 8'd202; b = 8'd239;  #10 
a = 8'd202; b = 8'd240;  #10 
a = 8'd202; b = 8'd241;  #10 
a = 8'd202; b = 8'd242;  #10 
a = 8'd202; b = 8'd243;  #10 
a = 8'd202; b = 8'd244;  #10 
a = 8'd202; b = 8'd245;  #10 
a = 8'd202; b = 8'd246;  #10 
a = 8'd202; b = 8'd247;  #10 
a = 8'd202; b = 8'd248;  #10 
a = 8'd202; b = 8'd249;  #10 
a = 8'd202; b = 8'd250;  #10 
a = 8'd202; b = 8'd251;  #10 
a = 8'd202; b = 8'd252;  #10 
a = 8'd202; b = 8'd253;  #10 
a = 8'd202; b = 8'd254;  #10 
a = 8'd202; b = 8'd255;  #10 
a = 8'd203; b = 8'd0;  #10 
a = 8'd203; b = 8'd1;  #10 
a = 8'd203; b = 8'd2;  #10 
a = 8'd203; b = 8'd3;  #10 
a = 8'd203; b = 8'd4;  #10 
a = 8'd203; b = 8'd5;  #10 
a = 8'd203; b = 8'd6;  #10 
a = 8'd203; b = 8'd7;  #10 
a = 8'd203; b = 8'd8;  #10 
a = 8'd203; b = 8'd9;  #10 
a = 8'd203; b = 8'd10;  #10 
a = 8'd203; b = 8'd11;  #10 
a = 8'd203; b = 8'd12;  #10 
a = 8'd203; b = 8'd13;  #10 
a = 8'd203; b = 8'd14;  #10 
a = 8'd203; b = 8'd15;  #10 
a = 8'd203; b = 8'd16;  #10 
a = 8'd203; b = 8'd17;  #10 
a = 8'd203; b = 8'd18;  #10 
a = 8'd203; b = 8'd19;  #10 
a = 8'd203; b = 8'd20;  #10 
a = 8'd203; b = 8'd21;  #10 
a = 8'd203; b = 8'd22;  #10 
a = 8'd203; b = 8'd23;  #10 
a = 8'd203; b = 8'd24;  #10 
a = 8'd203; b = 8'd25;  #10 
a = 8'd203; b = 8'd26;  #10 
a = 8'd203; b = 8'd27;  #10 
a = 8'd203; b = 8'd28;  #10 
a = 8'd203; b = 8'd29;  #10 
a = 8'd203; b = 8'd30;  #10 
a = 8'd203; b = 8'd31;  #10 
a = 8'd203; b = 8'd32;  #10 
a = 8'd203; b = 8'd33;  #10 
a = 8'd203; b = 8'd34;  #10 
a = 8'd203; b = 8'd35;  #10 
a = 8'd203; b = 8'd36;  #10 
a = 8'd203; b = 8'd37;  #10 
a = 8'd203; b = 8'd38;  #10 
a = 8'd203; b = 8'd39;  #10 
a = 8'd203; b = 8'd40;  #10 
a = 8'd203; b = 8'd41;  #10 
a = 8'd203; b = 8'd42;  #10 
a = 8'd203; b = 8'd43;  #10 
a = 8'd203; b = 8'd44;  #10 
a = 8'd203; b = 8'd45;  #10 
a = 8'd203; b = 8'd46;  #10 
a = 8'd203; b = 8'd47;  #10 
a = 8'd203; b = 8'd48;  #10 
a = 8'd203; b = 8'd49;  #10 
a = 8'd203; b = 8'd50;  #10 
a = 8'd203; b = 8'd51;  #10 
a = 8'd203; b = 8'd52;  #10 
a = 8'd203; b = 8'd53;  #10 
a = 8'd203; b = 8'd54;  #10 
a = 8'd203; b = 8'd55;  #10 
a = 8'd203; b = 8'd56;  #10 
a = 8'd203; b = 8'd57;  #10 
a = 8'd203; b = 8'd58;  #10 
a = 8'd203; b = 8'd59;  #10 
a = 8'd203; b = 8'd60;  #10 
a = 8'd203; b = 8'd61;  #10 
a = 8'd203; b = 8'd62;  #10 
a = 8'd203; b = 8'd63;  #10 
a = 8'd203; b = 8'd64;  #10 
a = 8'd203; b = 8'd65;  #10 
a = 8'd203; b = 8'd66;  #10 
a = 8'd203; b = 8'd67;  #10 
a = 8'd203; b = 8'd68;  #10 
a = 8'd203; b = 8'd69;  #10 
a = 8'd203; b = 8'd70;  #10 
a = 8'd203; b = 8'd71;  #10 
a = 8'd203; b = 8'd72;  #10 
a = 8'd203; b = 8'd73;  #10 
a = 8'd203; b = 8'd74;  #10 
a = 8'd203; b = 8'd75;  #10 
a = 8'd203; b = 8'd76;  #10 
a = 8'd203; b = 8'd77;  #10 
a = 8'd203; b = 8'd78;  #10 
a = 8'd203; b = 8'd79;  #10 
a = 8'd203; b = 8'd80;  #10 
a = 8'd203; b = 8'd81;  #10 
a = 8'd203; b = 8'd82;  #10 
a = 8'd203; b = 8'd83;  #10 
a = 8'd203; b = 8'd84;  #10 
a = 8'd203; b = 8'd85;  #10 
a = 8'd203; b = 8'd86;  #10 
a = 8'd203; b = 8'd87;  #10 
a = 8'd203; b = 8'd88;  #10 
a = 8'd203; b = 8'd89;  #10 
a = 8'd203; b = 8'd90;  #10 
a = 8'd203; b = 8'd91;  #10 
a = 8'd203; b = 8'd92;  #10 
a = 8'd203; b = 8'd93;  #10 
a = 8'd203; b = 8'd94;  #10 
a = 8'd203; b = 8'd95;  #10 
a = 8'd203; b = 8'd96;  #10 
a = 8'd203; b = 8'd97;  #10 
a = 8'd203; b = 8'd98;  #10 
a = 8'd203; b = 8'd99;  #10 
a = 8'd203; b = 8'd100;  #10 
a = 8'd203; b = 8'd101;  #10 
a = 8'd203; b = 8'd102;  #10 
a = 8'd203; b = 8'd103;  #10 
a = 8'd203; b = 8'd104;  #10 
a = 8'd203; b = 8'd105;  #10 
a = 8'd203; b = 8'd106;  #10 
a = 8'd203; b = 8'd107;  #10 
a = 8'd203; b = 8'd108;  #10 
a = 8'd203; b = 8'd109;  #10 
a = 8'd203; b = 8'd110;  #10 
a = 8'd203; b = 8'd111;  #10 
a = 8'd203; b = 8'd112;  #10 
a = 8'd203; b = 8'd113;  #10 
a = 8'd203; b = 8'd114;  #10 
a = 8'd203; b = 8'd115;  #10 
a = 8'd203; b = 8'd116;  #10 
a = 8'd203; b = 8'd117;  #10 
a = 8'd203; b = 8'd118;  #10 
a = 8'd203; b = 8'd119;  #10 
a = 8'd203; b = 8'd120;  #10 
a = 8'd203; b = 8'd121;  #10 
a = 8'd203; b = 8'd122;  #10 
a = 8'd203; b = 8'd123;  #10 
a = 8'd203; b = 8'd124;  #10 
a = 8'd203; b = 8'd125;  #10 
a = 8'd203; b = 8'd126;  #10 
a = 8'd203; b = 8'd127;  #10 
a = 8'd203; b = 8'd128;  #10 
a = 8'd203; b = 8'd129;  #10 
a = 8'd203; b = 8'd130;  #10 
a = 8'd203; b = 8'd131;  #10 
a = 8'd203; b = 8'd132;  #10 
a = 8'd203; b = 8'd133;  #10 
a = 8'd203; b = 8'd134;  #10 
a = 8'd203; b = 8'd135;  #10 
a = 8'd203; b = 8'd136;  #10 
a = 8'd203; b = 8'd137;  #10 
a = 8'd203; b = 8'd138;  #10 
a = 8'd203; b = 8'd139;  #10 
a = 8'd203; b = 8'd140;  #10 
a = 8'd203; b = 8'd141;  #10 
a = 8'd203; b = 8'd142;  #10 
a = 8'd203; b = 8'd143;  #10 
a = 8'd203; b = 8'd144;  #10 
a = 8'd203; b = 8'd145;  #10 
a = 8'd203; b = 8'd146;  #10 
a = 8'd203; b = 8'd147;  #10 
a = 8'd203; b = 8'd148;  #10 
a = 8'd203; b = 8'd149;  #10 
a = 8'd203; b = 8'd150;  #10 
a = 8'd203; b = 8'd151;  #10 
a = 8'd203; b = 8'd152;  #10 
a = 8'd203; b = 8'd153;  #10 
a = 8'd203; b = 8'd154;  #10 
a = 8'd203; b = 8'd155;  #10 
a = 8'd203; b = 8'd156;  #10 
a = 8'd203; b = 8'd157;  #10 
a = 8'd203; b = 8'd158;  #10 
a = 8'd203; b = 8'd159;  #10 
a = 8'd203; b = 8'd160;  #10 
a = 8'd203; b = 8'd161;  #10 
a = 8'd203; b = 8'd162;  #10 
a = 8'd203; b = 8'd163;  #10 
a = 8'd203; b = 8'd164;  #10 
a = 8'd203; b = 8'd165;  #10 
a = 8'd203; b = 8'd166;  #10 
a = 8'd203; b = 8'd167;  #10 
a = 8'd203; b = 8'd168;  #10 
a = 8'd203; b = 8'd169;  #10 
a = 8'd203; b = 8'd170;  #10 
a = 8'd203; b = 8'd171;  #10 
a = 8'd203; b = 8'd172;  #10 
a = 8'd203; b = 8'd173;  #10 
a = 8'd203; b = 8'd174;  #10 
a = 8'd203; b = 8'd175;  #10 
a = 8'd203; b = 8'd176;  #10 
a = 8'd203; b = 8'd177;  #10 
a = 8'd203; b = 8'd178;  #10 
a = 8'd203; b = 8'd179;  #10 
a = 8'd203; b = 8'd180;  #10 
a = 8'd203; b = 8'd181;  #10 
a = 8'd203; b = 8'd182;  #10 
a = 8'd203; b = 8'd183;  #10 
a = 8'd203; b = 8'd184;  #10 
a = 8'd203; b = 8'd185;  #10 
a = 8'd203; b = 8'd186;  #10 
a = 8'd203; b = 8'd187;  #10 
a = 8'd203; b = 8'd188;  #10 
a = 8'd203; b = 8'd189;  #10 
a = 8'd203; b = 8'd190;  #10 
a = 8'd203; b = 8'd191;  #10 
a = 8'd203; b = 8'd192;  #10 
a = 8'd203; b = 8'd193;  #10 
a = 8'd203; b = 8'd194;  #10 
a = 8'd203; b = 8'd195;  #10 
a = 8'd203; b = 8'd196;  #10 
a = 8'd203; b = 8'd197;  #10 
a = 8'd203; b = 8'd198;  #10 
a = 8'd203; b = 8'd199;  #10 
a = 8'd203; b = 8'd200;  #10 
a = 8'd203; b = 8'd201;  #10 
a = 8'd203; b = 8'd202;  #10 
a = 8'd203; b = 8'd203;  #10 
a = 8'd203; b = 8'd204;  #10 
a = 8'd203; b = 8'd205;  #10 
a = 8'd203; b = 8'd206;  #10 
a = 8'd203; b = 8'd207;  #10 
a = 8'd203; b = 8'd208;  #10 
a = 8'd203; b = 8'd209;  #10 
a = 8'd203; b = 8'd210;  #10 
a = 8'd203; b = 8'd211;  #10 
a = 8'd203; b = 8'd212;  #10 
a = 8'd203; b = 8'd213;  #10 
a = 8'd203; b = 8'd214;  #10 
a = 8'd203; b = 8'd215;  #10 
a = 8'd203; b = 8'd216;  #10 
a = 8'd203; b = 8'd217;  #10 
a = 8'd203; b = 8'd218;  #10 
a = 8'd203; b = 8'd219;  #10 
a = 8'd203; b = 8'd220;  #10 
a = 8'd203; b = 8'd221;  #10 
a = 8'd203; b = 8'd222;  #10 
a = 8'd203; b = 8'd223;  #10 
a = 8'd203; b = 8'd224;  #10 
a = 8'd203; b = 8'd225;  #10 
a = 8'd203; b = 8'd226;  #10 
a = 8'd203; b = 8'd227;  #10 
a = 8'd203; b = 8'd228;  #10 
a = 8'd203; b = 8'd229;  #10 
a = 8'd203; b = 8'd230;  #10 
a = 8'd203; b = 8'd231;  #10 
a = 8'd203; b = 8'd232;  #10 
a = 8'd203; b = 8'd233;  #10 
a = 8'd203; b = 8'd234;  #10 
a = 8'd203; b = 8'd235;  #10 
a = 8'd203; b = 8'd236;  #10 
a = 8'd203; b = 8'd237;  #10 
a = 8'd203; b = 8'd238;  #10 
a = 8'd203; b = 8'd239;  #10 
a = 8'd203; b = 8'd240;  #10 
a = 8'd203; b = 8'd241;  #10 
a = 8'd203; b = 8'd242;  #10 
a = 8'd203; b = 8'd243;  #10 
a = 8'd203; b = 8'd244;  #10 
a = 8'd203; b = 8'd245;  #10 
a = 8'd203; b = 8'd246;  #10 
a = 8'd203; b = 8'd247;  #10 
a = 8'd203; b = 8'd248;  #10 
a = 8'd203; b = 8'd249;  #10 
a = 8'd203; b = 8'd250;  #10 
a = 8'd203; b = 8'd251;  #10 
a = 8'd203; b = 8'd252;  #10 
a = 8'd203; b = 8'd253;  #10 
a = 8'd203; b = 8'd254;  #10 
a = 8'd203; b = 8'd255;  #10 
a = 8'd204; b = 8'd0;  #10 
a = 8'd204; b = 8'd1;  #10 
a = 8'd204; b = 8'd2;  #10 
a = 8'd204; b = 8'd3;  #10 
a = 8'd204; b = 8'd4;  #10 
a = 8'd204; b = 8'd5;  #10 
a = 8'd204; b = 8'd6;  #10 
a = 8'd204; b = 8'd7;  #10 
a = 8'd204; b = 8'd8;  #10 
a = 8'd204; b = 8'd9;  #10 
a = 8'd204; b = 8'd10;  #10 
a = 8'd204; b = 8'd11;  #10 
a = 8'd204; b = 8'd12;  #10 
a = 8'd204; b = 8'd13;  #10 
a = 8'd204; b = 8'd14;  #10 
a = 8'd204; b = 8'd15;  #10 
a = 8'd204; b = 8'd16;  #10 
a = 8'd204; b = 8'd17;  #10 
a = 8'd204; b = 8'd18;  #10 
a = 8'd204; b = 8'd19;  #10 
a = 8'd204; b = 8'd20;  #10 
a = 8'd204; b = 8'd21;  #10 
a = 8'd204; b = 8'd22;  #10 
a = 8'd204; b = 8'd23;  #10 
a = 8'd204; b = 8'd24;  #10 
a = 8'd204; b = 8'd25;  #10 
a = 8'd204; b = 8'd26;  #10 
a = 8'd204; b = 8'd27;  #10 
a = 8'd204; b = 8'd28;  #10 
a = 8'd204; b = 8'd29;  #10 
a = 8'd204; b = 8'd30;  #10 
a = 8'd204; b = 8'd31;  #10 
a = 8'd204; b = 8'd32;  #10 
a = 8'd204; b = 8'd33;  #10 
a = 8'd204; b = 8'd34;  #10 
a = 8'd204; b = 8'd35;  #10 
a = 8'd204; b = 8'd36;  #10 
a = 8'd204; b = 8'd37;  #10 
a = 8'd204; b = 8'd38;  #10 
a = 8'd204; b = 8'd39;  #10 
a = 8'd204; b = 8'd40;  #10 
a = 8'd204; b = 8'd41;  #10 
a = 8'd204; b = 8'd42;  #10 
a = 8'd204; b = 8'd43;  #10 
a = 8'd204; b = 8'd44;  #10 
a = 8'd204; b = 8'd45;  #10 
a = 8'd204; b = 8'd46;  #10 
a = 8'd204; b = 8'd47;  #10 
a = 8'd204; b = 8'd48;  #10 
a = 8'd204; b = 8'd49;  #10 
a = 8'd204; b = 8'd50;  #10 
a = 8'd204; b = 8'd51;  #10 
a = 8'd204; b = 8'd52;  #10 
a = 8'd204; b = 8'd53;  #10 
a = 8'd204; b = 8'd54;  #10 
a = 8'd204; b = 8'd55;  #10 
a = 8'd204; b = 8'd56;  #10 
a = 8'd204; b = 8'd57;  #10 
a = 8'd204; b = 8'd58;  #10 
a = 8'd204; b = 8'd59;  #10 
a = 8'd204; b = 8'd60;  #10 
a = 8'd204; b = 8'd61;  #10 
a = 8'd204; b = 8'd62;  #10 
a = 8'd204; b = 8'd63;  #10 
a = 8'd204; b = 8'd64;  #10 
a = 8'd204; b = 8'd65;  #10 
a = 8'd204; b = 8'd66;  #10 
a = 8'd204; b = 8'd67;  #10 
a = 8'd204; b = 8'd68;  #10 
a = 8'd204; b = 8'd69;  #10 
a = 8'd204; b = 8'd70;  #10 
a = 8'd204; b = 8'd71;  #10 
a = 8'd204; b = 8'd72;  #10 
a = 8'd204; b = 8'd73;  #10 
a = 8'd204; b = 8'd74;  #10 
a = 8'd204; b = 8'd75;  #10 
a = 8'd204; b = 8'd76;  #10 
a = 8'd204; b = 8'd77;  #10 
a = 8'd204; b = 8'd78;  #10 
a = 8'd204; b = 8'd79;  #10 
a = 8'd204; b = 8'd80;  #10 
a = 8'd204; b = 8'd81;  #10 
a = 8'd204; b = 8'd82;  #10 
a = 8'd204; b = 8'd83;  #10 
a = 8'd204; b = 8'd84;  #10 
a = 8'd204; b = 8'd85;  #10 
a = 8'd204; b = 8'd86;  #10 
a = 8'd204; b = 8'd87;  #10 
a = 8'd204; b = 8'd88;  #10 
a = 8'd204; b = 8'd89;  #10 
a = 8'd204; b = 8'd90;  #10 
a = 8'd204; b = 8'd91;  #10 
a = 8'd204; b = 8'd92;  #10 
a = 8'd204; b = 8'd93;  #10 
a = 8'd204; b = 8'd94;  #10 
a = 8'd204; b = 8'd95;  #10 
a = 8'd204; b = 8'd96;  #10 
a = 8'd204; b = 8'd97;  #10 
a = 8'd204; b = 8'd98;  #10 
a = 8'd204; b = 8'd99;  #10 
a = 8'd204; b = 8'd100;  #10 
a = 8'd204; b = 8'd101;  #10 
a = 8'd204; b = 8'd102;  #10 
a = 8'd204; b = 8'd103;  #10 
a = 8'd204; b = 8'd104;  #10 
a = 8'd204; b = 8'd105;  #10 
a = 8'd204; b = 8'd106;  #10 
a = 8'd204; b = 8'd107;  #10 
a = 8'd204; b = 8'd108;  #10 
a = 8'd204; b = 8'd109;  #10 
a = 8'd204; b = 8'd110;  #10 
a = 8'd204; b = 8'd111;  #10 
a = 8'd204; b = 8'd112;  #10 
a = 8'd204; b = 8'd113;  #10 
a = 8'd204; b = 8'd114;  #10 
a = 8'd204; b = 8'd115;  #10 
a = 8'd204; b = 8'd116;  #10 
a = 8'd204; b = 8'd117;  #10 
a = 8'd204; b = 8'd118;  #10 
a = 8'd204; b = 8'd119;  #10 
a = 8'd204; b = 8'd120;  #10 
a = 8'd204; b = 8'd121;  #10 
a = 8'd204; b = 8'd122;  #10 
a = 8'd204; b = 8'd123;  #10 
a = 8'd204; b = 8'd124;  #10 
a = 8'd204; b = 8'd125;  #10 
a = 8'd204; b = 8'd126;  #10 
a = 8'd204; b = 8'd127;  #10 
a = 8'd204; b = 8'd128;  #10 
a = 8'd204; b = 8'd129;  #10 
a = 8'd204; b = 8'd130;  #10 
a = 8'd204; b = 8'd131;  #10 
a = 8'd204; b = 8'd132;  #10 
a = 8'd204; b = 8'd133;  #10 
a = 8'd204; b = 8'd134;  #10 
a = 8'd204; b = 8'd135;  #10 
a = 8'd204; b = 8'd136;  #10 
a = 8'd204; b = 8'd137;  #10 
a = 8'd204; b = 8'd138;  #10 
a = 8'd204; b = 8'd139;  #10 
a = 8'd204; b = 8'd140;  #10 
a = 8'd204; b = 8'd141;  #10 
a = 8'd204; b = 8'd142;  #10 
a = 8'd204; b = 8'd143;  #10 
a = 8'd204; b = 8'd144;  #10 
a = 8'd204; b = 8'd145;  #10 
a = 8'd204; b = 8'd146;  #10 
a = 8'd204; b = 8'd147;  #10 
a = 8'd204; b = 8'd148;  #10 
a = 8'd204; b = 8'd149;  #10 
a = 8'd204; b = 8'd150;  #10 
a = 8'd204; b = 8'd151;  #10 
a = 8'd204; b = 8'd152;  #10 
a = 8'd204; b = 8'd153;  #10 
a = 8'd204; b = 8'd154;  #10 
a = 8'd204; b = 8'd155;  #10 
a = 8'd204; b = 8'd156;  #10 
a = 8'd204; b = 8'd157;  #10 
a = 8'd204; b = 8'd158;  #10 
a = 8'd204; b = 8'd159;  #10 
a = 8'd204; b = 8'd160;  #10 
a = 8'd204; b = 8'd161;  #10 
a = 8'd204; b = 8'd162;  #10 
a = 8'd204; b = 8'd163;  #10 
a = 8'd204; b = 8'd164;  #10 
a = 8'd204; b = 8'd165;  #10 
a = 8'd204; b = 8'd166;  #10 
a = 8'd204; b = 8'd167;  #10 
a = 8'd204; b = 8'd168;  #10 
a = 8'd204; b = 8'd169;  #10 
a = 8'd204; b = 8'd170;  #10 
a = 8'd204; b = 8'd171;  #10 
a = 8'd204; b = 8'd172;  #10 
a = 8'd204; b = 8'd173;  #10 
a = 8'd204; b = 8'd174;  #10 
a = 8'd204; b = 8'd175;  #10 
a = 8'd204; b = 8'd176;  #10 
a = 8'd204; b = 8'd177;  #10 
a = 8'd204; b = 8'd178;  #10 
a = 8'd204; b = 8'd179;  #10 
a = 8'd204; b = 8'd180;  #10 
a = 8'd204; b = 8'd181;  #10 
a = 8'd204; b = 8'd182;  #10 
a = 8'd204; b = 8'd183;  #10 
a = 8'd204; b = 8'd184;  #10 
a = 8'd204; b = 8'd185;  #10 
a = 8'd204; b = 8'd186;  #10 
a = 8'd204; b = 8'd187;  #10 
a = 8'd204; b = 8'd188;  #10 
a = 8'd204; b = 8'd189;  #10 
a = 8'd204; b = 8'd190;  #10 
a = 8'd204; b = 8'd191;  #10 
a = 8'd204; b = 8'd192;  #10 
a = 8'd204; b = 8'd193;  #10 
a = 8'd204; b = 8'd194;  #10 
a = 8'd204; b = 8'd195;  #10 
a = 8'd204; b = 8'd196;  #10 
a = 8'd204; b = 8'd197;  #10 
a = 8'd204; b = 8'd198;  #10 
a = 8'd204; b = 8'd199;  #10 
a = 8'd204; b = 8'd200;  #10 
a = 8'd204; b = 8'd201;  #10 
a = 8'd204; b = 8'd202;  #10 
a = 8'd204; b = 8'd203;  #10 
a = 8'd204; b = 8'd204;  #10 
a = 8'd204; b = 8'd205;  #10 
a = 8'd204; b = 8'd206;  #10 
a = 8'd204; b = 8'd207;  #10 
a = 8'd204; b = 8'd208;  #10 
a = 8'd204; b = 8'd209;  #10 
a = 8'd204; b = 8'd210;  #10 
a = 8'd204; b = 8'd211;  #10 
a = 8'd204; b = 8'd212;  #10 
a = 8'd204; b = 8'd213;  #10 
a = 8'd204; b = 8'd214;  #10 
a = 8'd204; b = 8'd215;  #10 
a = 8'd204; b = 8'd216;  #10 
a = 8'd204; b = 8'd217;  #10 
a = 8'd204; b = 8'd218;  #10 
a = 8'd204; b = 8'd219;  #10 
a = 8'd204; b = 8'd220;  #10 
a = 8'd204; b = 8'd221;  #10 
a = 8'd204; b = 8'd222;  #10 
a = 8'd204; b = 8'd223;  #10 
a = 8'd204; b = 8'd224;  #10 
a = 8'd204; b = 8'd225;  #10 
a = 8'd204; b = 8'd226;  #10 
a = 8'd204; b = 8'd227;  #10 
a = 8'd204; b = 8'd228;  #10 
a = 8'd204; b = 8'd229;  #10 
a = 8'd204; b = 8'd230;  #10 
a = 8'd204; b = 8'd231;  #10 
a = 8'd204; b = 8'd232;  #10 
a = 8'd204; b = 8'd233;  #10 
a = 8'd204; b = 8'd234;  #10 
a = 8'd204; b = 8'd235;  #10 
a = 8'd204; b = 8'd236;  #10 
a = 8'd204; b = 8'd237;  #10 
a = 8'd204; b = 8'd238;  #10 
a = 8'd204; b = 8'd239;  #10 
a = 8'd204; b = 8'd240;  #10 
a = 8'd204; b = 8'd241;  #10 
a = 8'd204; b = 8'd242;  #10 
a = 8'd204; b = 8'd243;  #10 
a = 8'd204; b = 8'd244;  #10 
a = 8'd204; b = 8'd245;  #10 
a = 8'd204; b = 8'd246;  #10 
a = 8'd204; b = 8'd247;  #10 
a = 8'd204; b = 8'd248;  #10 
a = 8'd204; b = 8'd249;  #10 
a = 8'd204; b = 8'd250;  #10 
a = 8'd204; b = 8'd251;  #10 
a = 8'd204; b = 8'd252;  #10 
a = 8'd204; b = 8'd253;  #10 
a = 8'd204; b = 8'd254;  #10 
a = 8'd204; b = 8'd255;  #10 
a = 8'd205; b = 8'd0;  #10 
a = 8'd205; b = 8'd1;  #10 
a = 8'd205; b = 8'd2;  #10 
a = 8'd205; b = 8'd3;  #10 
a = 8'd205; b = 8'd4;  #10 
a = 8'd205; b = 8'd5;  #10 
a = 8'd205; b = 8'd6;  #10 
a = 8'd205; b = 8'd7;  #10 
a = 8'd205; b = 8'd8;  #10 
a = 8'd205; b = 8'd9;  #10 
a = 8'd205; b = 8'd10;  #10 
a = 8'd205; b = 8'd11;  #10 
a = 8'd205; b = 8'd12;  #10 
a = 8'd205; b = 8'd13;  #10 
a = 8'd205; b = 8'd14;  #10 
a = 8'd205; b = 8'd15;  #10 
a = 8'd205; b = 8'd16;  #10 
a = 8'd205; b = 8'd17;  #10 
a = 8'd205; b = 8'd18;  #10 
a = 8'd205; b = 8'd19;  #10 
a = 8'd205; b = 8'd20;  #10 
a = 8'd205; b = 8'd21;  #10 
a = 8'd205; b = 8'd22;  #10 
a = 8'd205; b = 8'd23;  #10 
a = 8'd205; b = 8'd24;  #10 
a = 8'd205; b = 8'd25;  #10 
a = 8'd205; b = 8'd26;  #10 
a = 8'd205; b = 8'd27;  #10 
a = 8'd205; b = 8'd28;  #10 
a = 8'd205; b = 8'd29;  #10 
a = 8'd205; b = 8'd30;  #10 
a = 8'd205; b = 8'd31;  #10 
a = 8'd205; b = 8'd32;  #10 
a = 8'd205; b = 8'd33;  #10 
a = 8'd205; b = 8'd34;  #10 
a = 8'd205; b = 8'd35;  #10 
a = 8'd205; b = 8'd36;  #10 
a = 8'd205; b = 8'd37;  #10 
a = 8'd205; b = 8'd38;  #10 
a = 8'd205; b = 8'd39;  #10 
a = 8'd205; b = 8'd40;  #10 
a = 8'd205; b = 8'd41;  #10 
a = 8'd205; b = 8'd42;  #10 
a = 8'd205; b = 8'd43;  #10 
a = 8'd205; b = 8'd44;  #10 
a = 8'd205; b = 8'd45;  #10 
a = 8'd205; b = 8'd46;  #10 
a = 8'd205; b = 8'd47;  #10 
a = 8'd205; b = 8'd48;  #10 
a = 8'd205; b = 8'd49;  #10 
a = 8'd205; b = 8'd50;  #10 
a = 8'd205; b = 8'd51;  #10 
a = 8'd205; b = 8'd52;  #10 
a = 8'd205; b = 8'd53;  #10 
a = 8'd205; b = 8'd54;  #10 
a = 8'd205; b = 8'd55;  #10 
a = 8'd205; b = 8'd56;  #10 
a = 8'd205; b = 8'd57;  #10 
a = 8'd205; b = 8'd58;  #10 
a = 8'd205; b = 8'd59;  #10 
a = 8'd205; b = 8'd60;  #10 
a = 8'd205; b = 8'd61;  #10 
a = 8'd205; b = 8'd62;  #10 
a = 8'd205; b = 8'd63;  #10 
a = 8'd205; b = 8'd64;  #10 
a = 8'd205; b = 8'd65;  #10 
a = 8'd205; b = 8'd66;  #10 
a = 8'd205; b = 8'd67;  #10 
a = 8'd205; b = 8'd68;  #10 
a = 8'd205; b = 8'd69;  #10 
a = 8'd205; b = 8'd70;  #10 
a = 8'd205; b = 8'd71;  #10 
a = 8'd205; b = 8'd72;  #10 
a = 8'd205; b = 8'd73;  #10 
a = 8'd205; b = 8'd74;  #10 
a = 8'd205; b = 8'd75;  #10 
a = 8'd205; b = 8'd76;  #10 
a = 8'd205; b = 8'd77;  #10 
a = 8'd205; b = 8'd78;  #10 
a = 8'd205; b = 8'd79;  #10 
a = 8'd205; b = 8'd80;  #10 
a = 8'd205; b = 8'd81;  #10 
a = 8'd205; b = 8'd82;  #10 
a = 8'd205; b = 8'd83;  #10 
a = 8'd205; b = 8'd84;  #10 
a = 8'd205; b = 8'd85;  #10 
a = 8'd205; b = 8'd86;  #10 
a = 8'd205; b = 8'd87;  #10 
a = 8'd205; b = 8'd88;  #10 
a = 8'd205; b = 8'd89;  #10 
a = 8'd205; b = 8'd90;  #10 
a = 8'd205; b = 8'd91;  #10 
a = 8'd205; b = 8'd92;  #10 
a = 8'd205; b = 8'd93;  #10 
a = 8'd205; b = 8'd94;  #10 
a = 8'd205; b = 8'd95;  #10 
a = 8'd205; b = 8'd96;  #10 
a = 8'd205; b = 8'd97;  #10 
a = 8'd205; b = 8'd98;  #10 
a = 8'd205; b = 8'd99;  #10 
a = 8'd205; b = 8'd100;  #10 
a = 8'd205; b = 8'd101;  #10 
a = 8'd205; b = 8'd102;  #10 
a = 8'd205; b = 8'd103;  #10 
a = 8'd205; b = 8'd104;  #10 
a = 8'd205; b = 8'd105;  #10 
a = 8'd205; b = 8'd106;  #10 
a = 8'd205; b = 8'd107;  #10 
a = 8'd205; b = 8'd108;  #10 
a = 8'd205; b = 8'd109;  #10 
a = 8'd205; b = 8'd110;  #10 
a = 8'd205; b = 8'd111;  #10 
a = 8'd205; b = 8'd112;  #10 
a = 8'd205; b = 8'd113;  #10 
a = 8'd205; b = 8'd114;  #10 
a = 8'd205; b = 8'd115;  #10 
a = 8'd205; b = 8'd116;  #10 
a = 8'd205; b = 8'd117;  #10 
a = 8'd205; b = 8'd118;  #10 
a = 8'd205; b = 8'd119;  #10 
a = 8'd205; b = 8'd120;  #10 
a = 8'd205; b = 8'd121;  #10 
a = 8'd205; b = 8'd122;  #10 
a = 8'd205; b = 8'd123;  #10 
a = 8'd205; b = 8'd124;  #10 
a = 8'd205; b = 8'd125;  #10 
a = 8'd205; b = 8'd126;  #10 
a = 8'd205; b = 8'd127;  #10 
a = 8'd205; b = 8'd128;  #10 
a = 8'd205; b = 8'd129;  #10 
a = 8'd205; b = 8'd130;  #10 
a = 8'd205; b = 8'd131;  #10 
a = 8'd205; b = 8'd132;  #10 
a = 8'd205; b = 8'd133;  #10 
a = 8'd205; b = 8'd134;  #10 
a = 8'd205; b = 8'd135;  #10 
a = 8'd205; b = 8'd136;  #10 
a = 8'd205; b = 8'd137;  #10 
a = 8'd205; b = 8'd138;  #10 
a = 8'd205; b = 8'd139;  #10 
a = 8'd205; b = 8'd140;  #10 
a = 8'd205; b = 8'd141;  #10 
a = 8'd205; b = 8'd142;  #10 
a = 8'd205; b = 8'd143;  #10 
a = 8'd205; b = 8'd144;  #10 
a = 8'd205; b = 8'd145;  #10 
a = 8'd205; b = 8'd146;  #10 
a = 8'd205; b = 8'd147;  #10 
a = 8'd205; b = 8'd148;  #10 
a = 8'd205; b = 8'd149;  #10 
a = 8'd205; b = 8'd150;  #10 
a = 8'd205; b = 8'd151;  #10 
a = 8'd205; b = 8'd152;  #10 
a = 8'd205; b = 8'd153;  #10 
a = 8'd205; b = 8'd154;  #10 
a = 8'd205; b = 8'd155;  #10 
a = 8'd205; b = 8'd156;  #10 
a = 8'd205; b = 8'd157;  #10 
a = 8'd205; b = 8'd158;  #10 
a = 8'd205; b = 8'd159;  #10 
a = 8'd205; b = 8'd160;  #10 
a = 8'd205; b = 8'd161;  #10 
a = 8'd205; b = 8'd162;  #10 
a = 8'd205; b = 8'd163;  #10 
a = 8'd205; b = 8'd164;  #10 
a = 8'd205; b = 8'd165;  #10 
a = 8'd205; b = 8'd166;  #10 
a = 8'd205; b = 8'd167;  #10 
a = 8'd205; b = 8'd168;  #10 
a = 8'd205; b = 8'd169;  #10 
a = 8'd205; b = 8'd170;  #10 
a = 8'd205; b = 8'd171;  #10 
a = 8'd205; b = 8'd172;  #10 
a = 8'd205; b = 8'd173;  #10 
a = 8'd205; b = 8'd174;  #10 
a = 8'd205; b = 8'd175;  #10 
a = 8'd205; b = 8'd176;  #10 
a = 8'd205; b = 8'd177;  #10 
a = 8'd205; b = 8'd178;  #10 
a = 8'd205; b = 8'd179;  #10 
a = 8'd205; b = 8'd180;  #10 
a = 8'd205; b = 8'd181;  #10 
a = 8'd205; b = 8'd182;  #10 
a = 8'd205; b = 8'd183;  #10 
a = 8'd205; b = 8'd184;  #10 
a = 8'd205; b = 8'd185;  #10 
a = 8'd205; b = 8'd186;  #10 
a = 8'd205; b = 8'd187;  #10 
a = 8'd205; b = 8'd188;  #10 
a = 8'd205; b = 8'd189;  #10 
a = 8'd205; b = 8'd190;  #10 
a = 8'd205; b = 8'd191;  #10 
a = 8'd205; b = 8'd192;  #10 
a = 8'd205; b = 8'd193;  #10 
a = 8'd205; b = 8'd194;  #10 
a = 8'd205; b = 8'd195;  #10 
a = 8'd205; b = 8'd196;  #10 
a = 8'd205; b = 8'd197;  #10 
a = 8'd205; b = 8'd198;  #10 
a = 8'd205; b = 8'd199;  #10 
a = 8'd205; b = 8'd200;  #10 
a = 8'd205; b = 8'd201;  #10 
a = 8'd205; b = 8'd202;  #10 
a = 8'd205; b = 8'd203;  #10 
a = 8'd205; b = 8'd204;  #10 
a = 8'd205; b = 8'd205;  #10 
a = 8'd205; b = 8'd206;  #10 
a = 8'd205; b = 8'd207;  #10 
a = 8'd205; b = 8'd208;  #10 
a = 8'd205; b = 8'd209;  #10 
a = 8'd205; b = 8'd210;  #10 
a = 8'd205; b = 8'd211;  #10 
a = 8'd205; b = 8'd212;  #10 
a = 8'd205; b = 8'd213;  #10 
a = 8'd205; b = 8'd214;  #10 
a = 8'd205; b = 8'd215;  #10 
a = 8'd205; b = 8'd216;  #10 
a = 8'd205; b = 8'd217;  #10 
a = 8'd205; b = 8'd218;  #10 
a = 8'd205; b = 8'd219;  #10 
a = 8'd205; b = 8'd220;  #10 
a = 8'd205; b = 8'd221;  #10 
a = 8'd205; b = 8'd222;  #10 
a = 8'd205; b = 8'd223;  #10 
a = 8'd205; b = 8'd224;  #10 
a = 8'd205; b = 8'd225;  #10 
a = 8'd205; b = 8'd226;  #10 
a = 8'd205; b = 8'd227;  #10 
a = 8'd205; b = 8'd228;  #10 
a = 8'd205; b = 8'd229;  #10 
a = 8'd205; b = 8'd230;  #10 
a = 8'd205; b = 8'd231;  #10 
a = 8'd205; b = 8'd232;  #10 
a = 8'd205; b = 8'd233;  #10 
a = 8'd205; b = 8'd234;  #10 
a = 8'd205; b = 8'd235;  #10 
a = 8'd205; b = 8'd236;  #10 
a = 8'd205; b = 8'd237;  #10 
a = 8'd205; b = 8'd238;  #10 
a = 8'd205; b = 8'd239;  #10 
a = 8'd205; b = 8'd240;  #10 
a = 8'd205; b = 8'd241;  #10 
a = 8'd205; b = 8'd242;  #10 
a = 8'd205; b = 8'd243;  #10 
a = 8'd205; b = 8'd244;  #10 
a = 8'd205; b = 8'd245;  #10 
a = 8'd205; b = 8'd246;  #10 
a = 8'd205; b = 8'd247;  #10 
a = 8'd205; b = 8'd248;  #10 
a = 8'd205; b = 8'd249;  #10 
a = 8'd205; b = 8'd250;  #10 
a = 8'd205; b = 8'd251;  #10 
a = 8'd205; b = 8'd252;  #10 
a = 8'd205; b = 8'd253;  #10 
a = 8'd205; b = 8'd254;  #10 
a = 8'd205; b = 8'd255;  #10 
a = 8'd206; b = 8'd0;  #10 
a = 8'd206; b = 8'd1;  #10 
a = 8'd206; b = 8'd2;  #10 
a = 8'd206; b = 8'd3;  #10 
a = 8'd206; b = 8'd4;  #10 
a = 8'd206; b = 8'd5;  #10 
a = 8'd206; b = 8'd6;  #10 
a = 8'd206; b = 8'd7;  #10 
a = 8'd206; b = 8'd8;  #10 
a = 8'd206; b = 8'd9;  #10 
a = 8'd206; b = 8'd10;  #10 
a = 8'd206; b = 8'd11;  #10 
a = 8'd206; b = 8'd12;  #10 
a = 8'd206; b = 8'd13;  #10 
a = 8'd206; b = 8'd14;  #10 
a = 8'd206; b = 8'd15;  #10 
a = 8'd206; b = 8'd16;  #10 
a = 8'd206; b = 8'd17;  #10 
a = 8'd206; b = 8'd18;  #10 
a = 8'd206; b = 8'd19;  #10 
a = 8'd206; b = 8'd20;  #10 
a = 8'd206; b = 8'd21;  #10 
a = 8'd206; b = 8'd22;  #10 
a = 8'd206; b = 8'd23;  #10 
a = 8'd206; b = 8'd24;  #10 
a = 8'd206; b = 8'd25;  #10 
a = 8'd206; b = 8'd26;  #10 
a = 8'd206; b = 8'd27;  #10 
a = 8'd206; b = 8'd28;  #10 
a = 8'd206; b = 8'd29;  #10 
a = 8'd206; b = 8'd30;  #10 
a = 8'd206; b = 8'd31;  #10 
a = 8'd206; b = 8'd32;  #10 
a = 8'd206; b = 8'd33;  #10 
a = 8'd206; b = 8'd34;  #10 
a = 8'd206; b = 8'd35;  #10 
a = 8'd206; b = 8'd36;  #10 
a = 8'd206; b = 8'd37;  #10 
a = 8'd206; b = 8'd38;  #10 
a = 8'd206; b = 8'd39;  #10 
a = 8'd206; b = 8'd40;  #10 
a = 8'd206; b = 8'd41;  #10 
a = 8'd206; b = 8'd42;  #10 
a = 8'd206; b = 8'd43;  #10 
a = 8'd206; b = 8'd44;  #10 
a = 8'd206; b = 8'd45;  #10 
a = 8'd206; b = 8'd46;  #10 
a = 8'd206; b = 8'd47;  #10 
a = 8'd206; b = 8'd48;  #10 
a = 8'd206; b = 8'd49;  #10 
a = 8'd206; b = 8'd50;  #10 
a = 8'd206; b = 8'd51;  #10 
a = 8'd206; b = 8'd52;  #10 
a = 8'd206; b = 8'd53;  #10 
a = 8'd206; b = 8'd54;  #10 
a = 8'd206; b = 8'd55;  #10 
a = 8'd206; b = 8'd56;  #10 
a = 8'd206; b = 8'd57;  #10 
a = 8'd206; b = 8'd58;  #10 
a = 8'd206; b = 8'd59;  #10 
a = 8'd206; b = 8'd60;  #10 
a = 8'd206; b = 8'd61;  #10 
a = 8'd206; b = 8'd62;  #10 
a = 8'd206; b = 8'd63;  #10 
a = 8'd206; b = 8'd64;  #10 
a = 8'd206; b = 8'd65;  #10 
a = 8'd206; b = 8'd66;  #10 
a = 8'd206; b = 8'd67;  #10 
a = 8'd206; b = 8'd68;  #10 
a = 8'd206; b = 8'd69;  #10 
a = 8'd206; b = 8'd70;  #10 
a = 8'd206; b = 8'd71;  #10 
a = 8'd206; b = 8'd72;  #10 
a = 8'd206; b = 8'd73;  #10 
a = 8'd206; b = 8'd74;  #10 
a = 8'd206; b = 8'd75;  #10 
a = 8'd206; b = 8'd76;  #10 
a = 8'd206; b = 8'd77;  #10 
a = 8'd206; b = 8'd78;  #10 
a = 8'd206; b = 8'd79;  #10 
a = 8'd206; b = 8'd80;  #10 
a = 8'd206; b = 8'd81;  #10 
a = 8'd206; b = 8'd82;  #10 
a = 8'd206; b = 8'd83;  #10 
a = 8'd206; b = 8'd84;  #10 
a = 8'd206; b = 8'd85;  #10 
a = 8'd206; b = 8'd86;  #10 
a = 8'd206; b = 8'd87;  #10 
a = 8'd206; b = 8'd88;  #10 
a = 8'd206; b = 8'd89;  #10 
a = 8'd206; b = 8'd90;  #10 
a = 8'd206; b = 8'd91;  #10 
a = 8'd206; b = 8'd92;  #10 
a = 8'd206; b = 8'd93;  #10 
a = 8'd206; b = 8'd94;  #10 
a = 8'd206; b = 8'd95;  #10 
a = 8'd206; b = 8'd96;  #10 
a = 8'd206; b = 8'd97;  #10 
a = 8'd206; b = 8'd98;  #10 
a = 8'd206; b = 8'd99;  #10 
a = 8'd206; b = 8'd100;  #10 
a = 8'd206; b = 8'd101;  #10 
a = 8'd206; b = 8'd102;  #10 
a = 8'd206; b = 8'd103;  #10 
a = 8'd206; b = 8'd104;  #10 
a = 8'd206; b = 8'd105;  #10 
a = 8'd206; b = 8'd106;  #10 
a = 8'd206; b = 8'd107;  #10 
a = 8'd206; b = 8'd108;  #10 
a = 8'd206; b = 8'd109;  #10 
a = 8'd206; b = 8'd110;  #10 
a = 8'd206; b = 8'd111;  #10 
a = 8'd206; b = 8'd112;  #10 
a = 8'd206; b = 8'd113;  #10 
a = 8'd206; b = 8'd114;  #10 
a = 8'd206; b = 8'd115;  #10 
a = 8'd206; b = 8'd116;  #10 
a = 8'd206; b = 8'd117;  #10 
a = 8'd206; b = 8'd118;  #10 
a = 8'd206; b = 8'd119;  #10 
a = 8'd206; b = 8'd120;  #10 
a = 8'd206; b = 8'd121;  #10 
a = 8'd206; b = 8'd122;  #10 
a = 8'd206; b = 8'd123;  #10 
a = 8'd206; b = 8'd124;  #10 
a = 8'd206; b = 8'd125;  #10 
a = 8'd206; b = 8'd126;  #10 
a = 8'd206; b = 8'd127;  #10 
a = 8'd206; b = 8'd128;  #10 
a = 8'd206; b = 8'd129;  #10 
a = 8'd206; b = 8'd130;  #10 
a = 8'd206; b = 8'd131;  #10 
a = 8'd206; b = 8'd132;  #10 
a = 8'd206; b = 8'd133;  #10 
a = 8'd206; b = 8'd134;  #10 
a = 8'd206; b = 8'd135;  #10 
a = 8'd206; b = 8'd136;  #10 
a = 8'd206; b = 8'd137;  #10 
a = 8'd206; b = 8'd138;  #10 
a = 8'd206; b = 8'd139;  #10 
a = 8'd206; b = 8'd140;  #10 
a = 8'd206; b = 8'd141;  #10 
a = 8'd206; b = 8'd142;  #10 
a = 8'd206; b = 8'd143;  #10 
a = 8'd206; b = 8'd144;  #10 
a = 8'd206; b = 8'd145;  #10 
a = 8'd206; b = 8'd146;  #10 
a = 8'd206; b = 8'd147;  #10 
a = 8'd206; b = 8'd148;  #10 
a = 8'd206; b = 8'd149;  #10 
a = 8'd206; b = 8'd150;  #10 
a = 8'd206; b = 8'd151;  #10 
a = 8'd206; b = 8'd152;  #10 
a = 8'd206; b = 8'd153;  #10 
a = 8'd206; b = 8'd154;  #10 
a = 8'd206; b = 8'd155;  #10 
a = 8'd206; b = 8'd156;  #10 
a = 8'd206; b = 8'd157;  #10 
a = 8'd206; b = 8'd158;  #10 
a = 8'd206; b = 8'd159;  #10 
a = 8'd206; b = 8'd160;  #10 
a = 8'd206; b = 8'd161;  #10 
a = 8'd206; b = 8'd162;  #10 
a = 8'd206; b = 8'd163;  #10 
a = 8'd206; b = 8'd164;  #10 
a = 8'd206; b = 8'd165;  #10 
a = 8'd206; b = 8'd166;  #10 
a = 8'd206; b = 8'd167;  #10 
a = 8'd206; b = 8'd168;  #10 
a = 8'd206; b = 8'd169;  #10 
a = 8'd206; b = 8'd170;  #10 
a = 8'd206; b = 8'd171;  #10 
a = 8'd206; b = 8'd172;  #10 
a = 8'd206; b = 8'd173;  #10 
a = 8'd206; b = 8'd174;  #10 
a = 8'd206; b = 8'd175;  #10 
a = 8'd206; b = 8'd176;  #10 
a = 8'd206; b = 8'd177;  #10 
a = 8'd206; b = 8'd178;  #10 
a = 8'd206; b = 8'd179;  #10 
a = 8'd206; b = 8'd180;  #10 
a = 8'd206; b = 8'd181;  #10 
a = 8'd206; b = 8'd182;  #10 
a = 8'd206; b = 8'd183;  #10 
a = 8'd206; b = 8'd184;  #10 
a = 8'd206; b = 8'd185;  #10 
a = 8'd206; b = 8'd186;  #10 
a = 8'd206; b = 8'd187;  #10 
a = 8'd206; b = 8'd188;  #10 
a = 8'd206; b = 8'd189;  #10 
a = 8'd206; b = 8'd190;  #10 
a = 8'd206; b = 8'd191;  #10 
a = 8'd206; b = 8'd192;  #10 
a = 8'd206; b = 8'd193;  #10 
a = 8'd206; b = 8'd194;  #10 
a = 8'd206; b = 8'd195;  #10 
a = 8'd206; b = 8'd196;  #10 
a = 8'd206; b = 8'd197;  #10 
a = 8'd206; b = 8'd198;  #10 
a = 8'd206; b = 8'd199;  #10 
a = 8'd206; b = 8'd200;  #10 
a = 8'd206; b = 8'd201;  #10 
a = 8'd206; b = 8'd202;  #10 
a = 8'd206; b = 8'd203;  #10 
a = 8'd206; b = 8'd204;  #10 
a = 8'd206; b = 8'd205;  #10 
a = 8'd206; b = 8'd206;  #10 
a = 8'd206; b = 8'd207;  #10 
a = 8'd206; b = 8'd208;  #10 
a = 8'd206; b = 8'd209;  #10 
a = 8'd206; b = 8'd210;  #10 
a = 8'd206; b = 8'd211;  #10 
a = 8'd206; b = 8'd212;  #10 
a = 8'd206; b = 8'd213;  #10 
a = 8'd206; b = 8'd214;  #10 
a = 8'd206; b = 8'd215;  #10 
a = 8'd206; b = 8'd216;  #10 
a = 8'd206; b = 8'd217;  #10 
a = 8'd206; b = 8'd218;  #10 
a = 8'd206; b = 8'd219;  #10 
a = 8'd206; b = 8'd220;  #10 
a = 8'd206; b = 8'd221;  #10 
a = 8'd206; b = 8'd222;  #10 
a = 8'd206; b = 8'd223;  #10 
a = 8'd206; b = 8'd224;  #10 
a = 8'd206; b = 8'd225;  #10 
a = 8'd206; b = 8'd226;  #10 
a = 8'd206; b = 8'd227;  #10 
a = 8'd206; b = 8'd228;  #10 
a = 8'd206; b = 8'd229;  #10 
a = 8'd206; b = 8'd230;  #10 
a = 8'd206; b = 8'd231;  #10 
a = 8'd206; b = 8'd232;  #10 
a = 8'd206; b = 8'd233;  #10 
a = 8'd206; b = 8'd234;  #10 
a = 8'd206; b = 8'd235;  #10 
a = 8'd206; b = 8'd236;  #10 
a = 8'd206; b = 8'd237;  #10 
a = 8'd206; b = 8'd238;  #10 
a = 8'd206; b = 8'd239;  #10 
a = 8'd206; b = 8'd240;  #10 
a = 8'd206; b = 8'd241;  #10 
a = 8'd206; b = 8'd242;  #10 
a = 8'd206; b = 8'd243;  #10 
a = 8'd206; b = 8'd244;  #10 
a = 8'd206; b = 8'd245;  #10 
a = 8'd206; b = 8'd246;  #10 
a = 8'd206; b = 8'd247;  #10 
a = 8'd206; b = 8'd248;  #10 
a = 8'd206; b = 8'd249;  #10 
a = 8'd206; b = 8'd250;  #10 
a = 8'd206; b = 8'd251;  #10 
a = 8'd206; b = 8'd252;  #10 
a = 8'd206; b = 8'd253;  #10 
a = 8'd206; b = 8'd254;  #10 
a = 8'd206; b = 8'd255;  #10 
a = 8'd207; b = 8'd0;  #10 
a = 8'd207; b = 8'd1;  #10 
a = 8'd207; b = 8'd2;  #10 
a = 8'd207; b = 8'd3;  #10 
a = 8'd207; b = 8'd4;  #10 
a = 8'd207; b = 8'd5;  #10 
a = 8'd207; b = 8'd6;  #10 
a = 8'd207; b = 8'd7;  #10 
a = 8'd207; b = 8'd8;  #10 
a = 8'd207; b = 8'd9;  #10 
a = 8'd207; b = 8'd10;  #10 
a = 8'd207; b = 8'd11;  #10 
a = 8'd207; b = 8'd12;  #10 
a = 8'd207; b = 8'd13;  #10 
a = 8'd207; b = 8'd14;  #10 
a = 8'd207; b = 8'd15;  #10 
a = 8'd207; b = 8'd16;  #10 
a = 8'd207; b = 8'd17;  #10 
a = 8'd207; b = 8'd18;  #10 
a = 8'd207; b = 8'd19;  #10 
a = 8'd207; b = 8'd20;  #10 
a = 8'd207; b = 8'd21;  #10 
a = 8'd207; b = 8'd22;  #10 
a = 8'd207; b = 8'd23;  #10 
a = 8'd207; b = 8'd24;  #10 
a = 8'd207; b = 8'd25;  #10 
a = 8'd207; b = 8'd26;  #10 
a = 8'd207; b = 8'd27;  #10 
a = 8'd207; b = 8'd28;  #10 
a = 8'd207; b = 8'd29;  #10 
a = 8'd207; b = 8'd30;  #10 
a = 8'd207; b = 8'd31;  #10 
a = 8'd207; b = 8'd32;  #10 
a = 8'd207; b = 8'd33;  #10 
a = 8'd207; b = 8'd34;  #10 
a = 8'd207; b = 8'd35;  #10 
a = 8'd207; b = 8'd36;  #10 
a = 8'd207; b = 8'd37;  #10 
a = 8'd207; b = 8'd38;  #10 
a = 8'd207; b = 8'd39;  #10 
a = 8'd207; b = 8'd40;  #10 
a = 8'd207; b = 8'd41;  #10 
a = 8'd207; b = 8'd42;  #10 
a = 8'd207; b = 8'd43;  #10 
a = 8'd207; b = 8'd44;  #10 
a = 8'd207; b = 8'd45;  #10 
a = 8'd207; b = 8'd46;  #10 
a = 8'd207; b = 8'd47;  #10 
a = 8'd207; b = 8'd48;  #10 
a = 8'd207; b = 8'd49;  #10 
a = 8'd207; b = 8'd50;  #10 
a = 8'd207; b = 8'd51;  #10 
a = 8'd207; b = 8'd52;  #10 
a = 8'd207; b = 8'd53;  #10 
a = 8'd207; b = 8'd54;  #10 
a = 8'd207; b = 8'd55;  #10 
a = 8'd207; b = 8'd56;  #10 
a = 8'd207; b = 8'd57;  #10 
a = 8'd207; b = 8'd58;  #10 
a = 8'd207; b = 8'd59;  #10 
a = 8'd207; b = 8'd60;  #10 
a = 8'd207; b = 8'd61;  #10 
a = 8'd207; b = 8'd62;  #10 
a = 8'd207; b = 8'd63;  #10 
a = 8'd207; b = 8'd64;  #10 
a = 8'd207; b = 8'd65;  #10 
a = 8'd207; b = 8'd66;  #10 
a = 8'd207; b = 8'd67;  #10 
a = 8'd207; b = 8'd68;  #10 
a = 8'd207; b = 8'd69;  #10 
a = 8'd207; b = 8'd70;  #10 
a = 8'd207; b = 8'd71;  #10 
a = 8'd207; b = 8'd72;  #10 
a = 8'd207; b = 8'd73;  #10 
a = 8'd207; b = 8'd74;  #10 
a = 8'd207; b = 8'd75;  #10 
a = 8'd207; b = 8'd76;  #10 
a = 8'd207; b = 8'd77;  #10 
a = 8'd207; b = 8'd78;  #10 
a = 8'd207; b = 8'd79;  #10 
a = 8'd207; b = 8'd80;  #10 
a = 8'd207; b = 8'd81;  #10 
a = 8'd207; b = 8'd82;  #10 
a = 8'd207; b = 8'd83;  #10 
a = 8'd207; b = 8'd84;  #10 
a = 8'd207; b = 8'd85;  #10 
a = 8'd207; b = 8'd86;  #10 
a = 8'd207; b = 8'd87;  #10 
a = 8'd207; b = 8'd88;  #10 
a = 8'd207; b = 8'd89;  #10 
a = 8'd207; b = 8'd90;  #10 
a = 8'd207; b = 8'd91;  #10 
a = 8'd207; b = 8'd92;  #10 
a = 8'd207; b = 8'd93;  #10 
a = 8'd207; b = 8'd94;  #10 
a = 8'd207; b = 8'd95;  #10 
a = 8'd207; b = 8'd96;  #10 
a = 8'd207; b = 8'd97;  #10 
a = 8'd207; b = 8'd98;  #10 
a = 8'd207; b = 8'd99;  #10 
a = 8'd207; b = 8'd100;  #10 
a = 8'd207; b = 8'd101;  #10 
a = 8'd207; b = 8'd102;  #10 
a = 8'd207; b = 8'd103;  #10 
a = 8'd207; b = 8'd104;  #10 
a = 8'd207; b = 8'd105;  #10 
a = 8'd207; b = 8'd106;  #10 
a = 8'd207; b = 8'd107;  #10 
a = 8'd207; b = 8'd108;  #10 
a = 8'd207; b = 8'd109;  #10 
a = 8'd207; b = 8'd110;  #10 
a = 8'd207; b = 8'd111;  #10 
a = 8'd207; b = 8'd112;  #10 
a = 8'd207; b = 8'd113;  #10 
a = 8'd207; b = 8'd114;  #10 
a = 8'd207; b = 8'd115;  #10 
a = 8'd207; b = 8'd116;  #10 
a = 8'd207; b = 8'd117;  #10 
a = 8'd207; b = 8'd118;  #10 
a = 8'd207; b = 8'd119;  #10 
a = 8'd207; b = 8'd120;  #10 
a = 8'd207; b = 8'd121;  #10 
a = 8'd207; b = 8'd122;  #10 
a = 8'd207; b = 8'd123;  #10 
a = 8'd207; b = 8'd124;  #10 
a = 8'd207; b = 8'd125;  #10 
a = 8'd207; b = 8'd126;  #10 
a = 8'd207; b = 8'd127;  #10 
a = 8'd207; b = 8'd128;  #10 
a = 8'd207; b = 8'd129;  #10 
a = 8'd207; b = 8'd130;  #10 
a = 8'd207; b = 8'd131;  #10 
a = 8'd207; b = 8'd132;  #10 
a = 8'd207; b = 8'd133;  #10 
a = 8'd207; b = 8'd134;  #10 
a = 8'd207; b = 8'd135;  #10 
a = 8'd207; b = 8'd136;  #10 
a = 8'd207; b = 8'd137;  #10 
a = 8'd207; b = 8'd138;  #10 
a = 8'd207; b = 8'd139;  #10 
a = 8'd207; b = 8'd140;  #10 
a = 8'd207; b = 8'd141;  #10 
a = 8'd207; b = 8'd142;  #10 
a = 8'd207; b = 8'd143;  #10 
a = 8'd207; b = 8'd144;  #10 
a = 8'd207; b = 8'd145;  #10 
a = 8'd207; b = 8'd146;  #10 
a = 8'd207; b = 8'd147;  #10 
a = 8'd207; b = 8'd148;  #10 
a = 8'd207; b = 8'd149;  #10 
a = 8'd207; b = 8'd150;  #10 
a = 8'd207; b = 8'd151;  #10 
a = 8'd207; b = 8'd152;  #10 
a = 8'd207; b = 8'd153;  #10 
a = 8'd207; b = 8'd154;  #10 
a = 8'd207; b = 8'd155;  #10 
a = 8'd207; b = 8'd156;  #10 
a = 8'd207; b = 8'd157;  #10 
a = 8'd207; b = 8'd158;  #10 
a = 8'd207; b = 8'd159;  #10 
a = 8'd207; b = 8'd160;  #10 
a = 8'd207; b = 8'd161;  #10 
a = 8'd207; b = 8'd162;  #10 
a = 8'd207; b = 8'd163;  #10 
a = 8'd207; b = 8'd164;  #10 
a = 8'd207; b = 8'd165;  #10 
a = 8'd207; b = 8'd166;  #10 
a = 8'd207; b = 8'd167;  #10 
a = 8'd207; b = 8'd168;  #10 
a = 8'd207; b = 8'd169;  #10 
a = 8'd207; b = 8'd170;  #10 
a = 8'd207; b = 8'd171;  #10 
a = 8'd207; b = 8'd172;  #10 
a = 8'd207; b = 8'd173;  #10 
a = 8'd207; b = 8'd174;  #10 
a = 8'd207; b = 8'd175;  #10 
a = 8'd207; b = 8'd176;  #10 
a = 8'd207; b = 8'd177;  #10 
a = 8'd207; b = 8'd178;  #10 
a = 8'd207; b = 8'd179;  #10 
a = 8'd207; b = 8'd180;  #10 
a = 8'd207; b = 8'd181;  #10 
a = 8'd207; b = 8'd182;  #10 
a = 8'd207; b = 8'd183;  #10 
a = 8'd207; b = 8'd184;  #10 
a = 8'd207; b = 8'd185;  #10 
a = 8'd207; b = 8'd186;  #10 
a = 8'd207; b = 8'd187;  #10 
a = 8'd207; b = 8'd188;  #10 
a = 8'd207; b = 8'd189;  #10 
a = 8'd207; b = 8'd190;  #10 
a = 8'd207; b = 8'd191;  #10 
a = 8'd207; b = 8'd192;  #10 
a = 8'd207; b = 8'd193;  #10 
a = 8'd207; b = 8'd194;  #10 
a = 8'd207; b = 8'd195;  #10 
a = 8'd207; b = 8'd196;  #10 
a = 8'd207; b = 8'd197;  #10 
a = 8'd207; b = 8'd198;  #10 
a = 8'd207; b = 8'd199;  #10 
a = 8'd207; b = 8'd200;  #10 
a = 8'd207; b = 8'd201;  #10 
a = 8'd207; b = 8'd202;  #10 
a = 8'd207; b = 8'd203;  #10 
a = 8'd207; b = 8'd204;  #10 
a = 8'd207; b = 8'd205;  #10 
a = 8'd207; b = 8'd206;  #10 
a = 8'd207; b = 8'd207;  #10 
a = 8'd207; b = 8'd208;  #10 
a = 8'd207; b = 8'd209;  #10 
a = 8'd207; b = 8'd210;  #10 
a = 8'd207; b = 8'd211;  #10 
a = 8'd207; b = 8'd212;  #10 
a = 8'd207; b = 8'd213;  #10 
a = 8'd207; b = 8'd214;  #10 
a = 8'd207; b = 8'd215;  #10 
a = 8'd207; b = 8'd216;  #10 
a = 8'd207; b = 8'd217;  #10 
a = 8'd207; b = 8'd218;  #10 
a = 8'd207; b = 8'd219;  #10 
a = 8'd207; b = 8'd220;  #10 
a = 8'd207; b = 8'd221;  #10 
a = 8'd207; b = 8'd222;  #10 
a = 8'd207; b = 8'd223;  #10 
a = 8'd207; b = 8'd224;  #10 
a = 8'd207; b = 8'd225;  #10 
a = 8'd207; b = 8'd226;  #10 
a = 8'd207; b = 8'd227;  #10 
a = 8'd207; b = 8'd228;  #10 
a = 8'd207; b = 8'd229;  #10 
a = 8'd207; b = 8'd230;  #10 
a = 8'd207; b = 8'd231;  #10 
a = 8'd207; b = 8'd232;  #10 
a = 8'd207; b = 8'd233;  #10 
a = 8'd207; b = 8'd234;  #10 
a = 8'd207; b = 8'd235;  #10 
a = 8'd207; b = 8'd236;  #10 
a = 8'd207; b = 8'd237;  #10 
a = 8'd207; b = 8'd238;  #10 
a = 8'd207; b = 8'd239;  #10 
a = 8'd207; b = 8'd240;  #10 
a = 8'd207; b = 8'd241;  #10 
a = 8'd207; b = 8'd242;  #10 
a = 8'd207; b = 8'd243;  #10 
a = 8'd207; b = 8'd244;  #10 
a = 8'd207; b = 8'd245;  #10 
a = 8'd207; b = 8'd246;  #10 
a = 8'd207; b = 8'd247;  #10 
a = 8'd207; b = 8'd248;  #10 
a = 8'd207; b = 8'd249;  #10 
a = 8'd207; b = 8'd250;  #10 
a = 8'd207; b = 8'd251;  #10 
a = 8'd207; b = 8'd252;  #10 
a = 8'd207; b = 8'd253;  #10 
a = 8'd207; b = 8'd254;  #10 
a = 8'd207; b = 8'd255;  #10 
a = 8'd208; b = 8'd0;  #10 
a = 8'd208; b = 8'd1;  #10 
a = 8'd208; b = 8'd2;  #10 
a = 8'd208; b = 8'd3;  #10 
a = 8'd208; b = 8'd4;  #10 
a = 8'd208; b = 8'd5;  #10 
a = 8'd208; b = 8'd6;  #10 
a = 8'd208; b = 8'd7;  #10 
a = 8'd208; b = 8'd8;  #10 
a = 8'd208; b = 8'd9;  #10 
a = 8'd208; b = 8'd10;  #10 
a = 8'd208; b = 8'd11;  #10 
a = 8'd208; b = 8'd12;  #10 
a = 8'd208; b = 8'd13;  #10 
a = 8'd208; b = 8'd14;  #10 
a = 8'd208; b = 8'd15;  #10 
a = 8'd208; b = 8'd16;  #10 
a = 8'd208; b = 8'd17;  #10 
a = 8'd208; b = 8'd18;  #10 
a = 8'd208; b = 8'd19;  #10 
a = 8'd208; b = 8'd20;  #10 
a = 8'd208; b = 8'd21;  #10 
a = 8'd208; b = 8'd22;  #10 
a = 8'd208; b = 8'd23;  #10 
a = 8'd208; b = 8'd24;  #10 
a = 8'd208; b = 8'd25;  #10 
a = 8'd208; b = 8'd26;  #10 
a = 8'd208; b = 8'd27;  #10 
a = 8'd208; b = 8'd28;  #10 
a = 8'd208; b = 8'd29;  #10 
a = 8'd208; b = 8'd30;  #10 
a = 8'd208; b = 8'd31;  #10 
a = 8'd208; b = 8'd32;  #10 
a = 8'd208; b = 8'd33;  #10 
a = 8'd208; b = 8'd34;  #10 
a = 8'd208; b = 8'd35;  #10 
a = 8'd208; b = 8'd36;  #10 
a = 8'd208; b = 8'd37;  #10 
a = 8'd208; b = 8'd38;  #10 
a = 8'd208; b = 8'd39;  #10 
a = 8'd208; b = 8'd40;  #10 
a = 8'd208; b = 8'd41;  #10 
a = 8'd208; b = 8'd42;  #10 
a = 8'd208; b = 8'd43;  #10 
a = 8'd208; b = 8'd44;  #10 
a = 8'd208; b = 8'd45;  #10 
a = 8'd208; b = 8'd46;  #10 
a = 8'd208; b = 8'd47;  #10 
a = 8'd208; b = 8'd48;  #10 
a = 8'd208; b = 8'd49;  #10 
a = 8'd208; b = 8'd50;  #10 
a = 8'd208; b = 8'd51;  #10 
a = 8'd208; b = 8'd52;  #10 
a = 8'd208; b = 8'd53;  #10 
a = 8'd208; b = 8'd54;  #10 
a = 8'd208; b = 8'd55;  #10 
a = 8'd208; b = 8'd56;  #10 
a = 8'd208; b = 8'd57;  #10 
a = 8'd208; b = 8'd58;  #10 
a = 8'd208; b = 8'd59;  #10 
a = 8'd208; b = 8'd60;  #10 
a = 8'd208; b = 8'd61;  #10 
a = 8'd208; b = 8'd62;  #10 
a = 8'd208; b = 8'd63;  #10 
a = 8'd208; b = 8'd64;  #10 
a = 8'd208; b = 8'd65;  #10 
a = 8'd208; b = 8'd66;  #10 
a = 8'd208; b = 8'd67;  #10 
a = 8'd208; b = 8'd68;  #10 
a = 8'd208; b = 8'd69;  #10 
a = 8'd208; b = 8'd70;  #10 
a = 8'd208; b = 8'd71;  #10 
a = 8'd208; b = 8'd72;  #10 
a = 8'd208; b = 8'd73;  #10 
a = 8'd208; b = 8'd74;  #10 
a = 8'd208; b = 8'd75;  #10 
a = 8'd208; b = 8'd76;  #10 
a = 8'd208; b = 8'd77;  #10 
a = 8'd208; b = 8'd78;  #10 
a = 8'd208; b = 8'd79;  #10 
a = 8'd208; b = 8'd80;  #10 
a = 8'd208; b = 8'd81;  #10 
a = 8'd208; b = 8'd82;  #10 
a = 8'd208; b = 8'd83;  #10 
a = 8'd208; b = 8'd84;  #10 
a = 8'd208; b = 8'd85;  #10 
a = 8'd208; b = 8'd86;  #10 
a = 8'd208; b = 8'd87;  #10 
a = 8'd208; b = 8'd88;  #10 
a = 8'd208; b = 8'd89;  #10 
a = 8'd208; b = 8'd90;  #10 
a = 8'd208; b = 8'd91;  #10 
a = 8'd208; b = 8'd92;  #10 
a = 8'd208; b = 8'd93;  #10 
a = 8'd208; b = 8'd94;  #10 
a = 8'd208; b = 8'd95;  #10 
a = 8'd208; b = 8'd96;  #10 
a = 8'd208; b = 8'd97;  #10 
a = 8'd208; b = 8'd98;  #10 
a = 8'd208; b = 8'd99;  #10 
a = 8'd208; b = 8'd100;  #10 
a = 8'd208; b = 8'd101;  #10 
a = 8'd208; b = 8'd102;  #10 
a = 8'd208; b = 8'd103;  #10 
a = 8'd208; b = 8'd104;  #10 
a = 8'd208; b = 8'd105;  #10 
a = 8'd208; b = 8'd106;  #10 
a = 8'd208; b = 8'd107;  #10 
a = 8'd208; b = 8'd108;  #10 
a = 8'd208; b = 8'd109;  #10 
a = 8'd208; b = 8'd110;  #10 
a = 8'd208; b = 8'd111;  #10 
a = 8'd208; b = 8'd112;  #10 
a = 8'd208; b = 8'd113;  #10 
a = 8'd208; b = 8'd114;  #10 
a = 8'd208; b = 8'd115;  #10 
a = 8'd208; b = 8'd116;  #10 
a = 8'd208; b = 8'd117;  #10 
a = 8'd208; b = 8'd118;  #10 
a = 8'd208; b = 8'd119;  #10 
a = 8'd208; b = 8'd120;  #10 
a = 8'd208; b = 8'd121;  #10 
a = 8'd208; b = 8'd122;  #10 
a = 8'd208; b = 8'd123;  #10 
a = 8'd208; b = 8'd124;  #10 
a = 8'd208; b = 8'd125;  #10 
a = 8'd208; b = 8'd126;  #10 
a = 8'd208; b = 8'd127;  #10 
a = 8'd208; b = 8'd128;  #10 
a = 8'd208; b = 8'd129;  #10 
a = 8'd208; b = 8'd130;  #10 
a = 8'd208; b = 8'd131;  #10 
a = 8'd208; b = 8'd132;  #10 
a = 8'd208; b = 8'd133;  #10 
a = 8'd208; b = 8'd134;  #10 
a = 8'd208; b = 8'd135;  #10 
a = 8'd208; b = 8'd136;  #10 
a = 8'd208; b = 8'd137;  #10 
a = 8'd208; b = 8'd138;  #10 
a = 8'd208; b = 8'd139;  #10 
a = 8'd208; b = 8'd140;  #10 
a = 8'd208; b = 8'd141;  #10 
a = 8'd208; b = 8'd142;  #10 
a = 8'd208; b = 8'd143;  #10 
a = 8'd208; b = 8'd144;  #10 
a = 8'd208; b = 8'd145;  #10 
a = 8'd208; b = 8'd146;  #10 
a = 8'd208; b = 8'd147;  #10 
a = 8'd208; b = 8'd148;  #10 
a = 8'd208; b = 8'd149;  #10 
a = 8'd208; b = 8'd150;  #10 
a = 8'd208; b = 8'd151;  #10 
a = 8'd208; b = 8'd152;  #10 
a = 8'd208; b = 8'd153;  #10 
a = 8'd208; b = 8'd154;  #10 
a = 8'd208; b = 8'd155;  #10 
a = 8'd208; b = 8'd156;  #10 
a = 8'd208; b = 8'd157;  #10 
a = 8'd208; b = 8'd158;  #10 
a = 8'd208; b = 8'd159;  #10 
a = 8'd208; b = 8'd160;  #10 
a = 8'd208; b = 8'd161;  #10 
a = 8'd208; b = 8'd162;  #10 
a = 8'd208; b = 8'd163;  #10 
a = 8'd208; b = 8'd164;  #10 
a = 8'd208; b = 8'd165;  #10 
a = 8'd208; b = 8'd166;  #10 
a = 8'd208; b = 8'd167;  #10 
a = 8'd208; b = 8'd168;  #10 
a = 8'd208; b = 8'd169;  #10 
a = 8'd208; b = 8'd170;  #10 
a = 8'd208; b = 8'd171;  #10 
a = 8'd208; b = 8'd172;  #10 
a = 8'd208; b = 8'd173;  #10 
a = 8'd208; b = 8'd174;  #10 
a = 8'd208; b = 8'd175;  #10 
a = 8'd208; b = 8'd176;  #10 
a = 8'd208; b = 8'd177;  #10 
a = 8'd208; b = 8'd178;  #10 
a = 8'd208; b = 8'd179;  #10 
a = 8'd208; b = 8'd180;  #10 
a = 8'd208; b = 8'd181;  #10 
a = 8'd208; b = 8'd182;  #10 
a = 8'd208; b = 8'd183;  #10 
a = 8'd208; b = 8'd184;  #10 
a = 8'd208; b = 8'd185;  #10 
a = 8'd208; b = 8'd186;  #10 
a = 8'd208; b = 8'd187;  #10 
a = 8'd208; b = 8'd188;  #10 
a = 8'd208; b = 8'd189;  #10 
a = 8'd208; b = 8'd190;  #10 
a = 8'd208; b = 8'd191;  #10 
a = 8'd208; b = 8'd192;  #10 
a = 8'd208; b = 8'd193;  #10 
a = 8'd208; b = 8'd194;  #10 
a = 8'd208; b = 8'd195;  #10 
a = 8'd208; b = 8'd196;  #10 
a = 8'd208; b = 8'd197;  #10 
a = 8'd208; b = 8'd198;  #10 
a = 8'd208; b = 8'd199;  #10 
a = 8'd208; b = 8'd200;  #10 
a = 8'd208; b = 8'd201;  #10 
a = 8'd208; b = 8'd202;  #10 
a = 8'd208; b = 8'd203;  #10 
a = 8'd208; b = 8'd204;  #10 
a = 8'd208; b = 8'd205;  #10 
a = 8'd208; b = 8'd206;  #10 
a = 8'd208; b = 8'd207;  #10 
a = 8'd208; b = 8'd208;  #10 
a = 8'd208; b = 8'd209;  #10 
a = 8'd208; b = 8'd210;  #10 
a = 8'd208; b = 8'd211;  #10 
a = 8'd208; b = 8'd212;  #10 
a = 8'd208; b = 8'd213;  #10 
a = 8'd208; b = 8'd214;  #10 
a = 8'd208; b = 8'd215;  #10 
a = 8'd208; b = 8'd216;  #10 
a = 8'd208; b = 8'd217;  #10 
a = 8'd208; b = 8'd218;  #10 
a = 8'd208; b = 8'd219;  #10 
a = 8'd208; b = 8'd220;  #10 
a = 8'd208; b = 8'd221;  #10 
a = 8'd208; b = 8'd222;  #10 
a = 8'd208; b = 8'd223;  #10 
a = 8'd208; b = 8'd224;  #10 
a = 8'd208; b = 8'd225;  #10 
a = 8'd208; b = 8'd226;  #10 
a = 8'd208; b = 8'd227;  #10 
a = 8'd208; b = 8'd228;  #10 
a = 8'd208; b = 8'd229;  #10 
a = 8'd208; b = 8'd230;  #10 
a = 8'd208; b = 8'd231;  #10 
a = 8'd208; b = 8'd232;  #10 
a = 8'd208; b = 8'd233;  #10 
a = 8'd208; b = 8'd234;  #10 
a = 8'd208; b = 8'd235;  #10 
a = 8'd208; b = 8'd236;  #10 
a = 8'd208; b = 8'd237;  #10 
a = 8'd208; b = 8'd238;  #10 
a = 8'd208; b = 8'd239;  #10 
a = 8'd208; b = 8'd240;  #10 
a = 8'd208; b = 8'd241;  #10 
a = 8'd208; b = 8'd242;  #10 
a = 8'd208; b = 8'd243;  #10 
a = 8'd208; b = 8'd244;  #10 
a = 8'd208; b = 8'd245;  #10 
a = 8'd208; b = 8'd246;  #10 
a = 8'd208; b = 8'd247;  #10 
a = 8'd208; b = 8'd248;  #10 
a = 8'd208; b = 8'd249;  #10 
a = 8'd208; b = 8'd250;  #10 
a = 8'd208; b = 8'd251;  #10 
a = 8'd208; b = 8'd252;  #10 
a = 8'd208; b = 8'd253;  #10 
a = 8'd208; b = 8'd254;  #10 
a = 8'd208; b = 8'd255;  #10 
a = 8'd209; b = 8'd0;  #10 
a = 8'd209; b = 8'd1;  #10 
a = 8'd209; b = 8'd2;  #10 
a = 8'd209; b = 8'd3;  #10 
a = 8'd209; b = 8'd4;  #10 
a = 8'd209; b = 8'd5;  #10 
a = 8'd209; b = 8'd6;  #10 
a = 8'd209; b = 8'd7;  #10 
a = 8'd209; b = 8'd8;  #10 
a = 8'd209; b = 8'd9;  #10 
a = 8'd209; b = 8'd10;  #10 
a = 8'd209; b = 8'd11;  #10 
a = 8'd209; b = 8'd12;  #10 
a = 8'd209; b = 8'd13;  #10 
a = 8'd209; b = 8'd14;  #10 
a = 8'd209; b = 8'd15;  #10 
a = 8'd209; b = 8'd16;  #10 
a = 8'd209; b = 8'd17;  #10 
a = 8'd209; b = 8'd18;  #10 
a = 8'd209; b = 8'd19;  #10 
a = 8'd209; b = 8'd20;  #10 
a = 8'd209; b = 8'd21;  #10 
a = 8'd209; b = 8'd22;  #10 
a = 8'd209; b = 8'd23;  #10 
a = 8'd209; b = 8'd24;  #10 
a = 8'd209; b = 8'd25;  #10 
a = 8'd209; b = 8'd26;  #10 
a = 8'd209; b = 8'd27;  #10 
a = 8'd209; b = 8'd28;  #10 
a = 8'd209; b = 8'd29;  #10 
a = 8'd209; b = 8'd30;  #10 
a = 8'd209; b = 8'd31;  #10 
a = 8'd209; b = 8'd32;  #10 
a = 8'd209; b = 8'd33;  #10 
a = 8'd209; b = 8'd34;  #10 
a = 8'd209; b = 8'd35;  #10 
a = 8'd209; b = 8'd36;  #10 
a = 8'd209; b = 8'd37;  #10 
a = 8'd209; b = 8'd38;  #10 
a = 8'd209; b = 8'd39;  #10 
a = 8'd209; b = 8'd40;  #10 
a = 8'd209; b = 8'd41;  #10 
a = 8'd209; b = 8'd42;  #10 
a = 8'd209; b = 8'd43;  #10 
a = 8'd209; b = 8'd44;  #10 
a = 8'd209; b = 8'd45;  #10 
a = 8'd209; b = 8'd46;  #10 
a = 8'd209; b = 8'd47;  #10 
a = 8'd209; b = 8'd48;  #10 
a = 8'd209; b = 8'd49;  #10 
a = 8'd209; b = 8'd50;  #10 
a = 8'd209; b = 8'd51;  #10 
a = 8'd209; b = 8'd52;  #10 
a = 8'd209; b = 8'd53;  #10 
a = 8'd209; b = 8'd54;  #10 
a = 8'd209; b = 8'd55;  #10 
a = 8'd209; b = 8'd56;  #10 
a = 8'd209; b = 8'd57;  #10 
a = 8'd209; b = 8'd58;  #10 
a = 8'd209; b = 8'd59;  #10 
a = 8'd209; b = 8'd60;  #10 
a = 8'd209; b = 8'd61;  #10 
a = 8'd209; b = 8'd62;  #10 
a = 8'd209; b = 8'd63;  #10 
a = 8'd209; b = 8'd64;  #10 
a = 8'd209; b = 8'd65;  #10 
a = 8'd209; b = 8'd66;  #10 
a = 8'd209; b = 8'd67;  #10 
a = 8'd209; b = 8'd68;  #10 
a = 8'd209; b = 8'd69;  #10 
a = 8'd209; b = 8'd70;  #10 
a = 8'd209; b = 8'd71;  #10 
a = 8'd209; b = 8'd72;  #10 
a = 8'd209; b = 8'd73;  #10 
a = 8'd209; b = 8'd74;  #10 
a = 8'd209; b = 8'd75;  #10 
a = 8'd209; b = 8'd76;  #10 
a = 8'd209; b = 8'd77;  #10 
a = 8'd209; b = 8'd78;  #10 
a = 8'd209; b = 8'd79;  #10 
a = 8'd209; b = 8'd80;  #10 
a = 8'd209; b = 8'd81;  #10 
a = 8'd209; b = 8'd82;  #10 
a = 8'd209; b = 8'd83;  #10 
a = 8'd209; b = 8'd84;  #10 
a = 8'd209; b = 8'd85;  #10 
a = 8'd209; b = 8'd86;  #10 
a = 8'd209; b = 8'd87;  #10 
a = 8'd209; b = 8'd88;  #10 
a = 8'd209; b = 8'd89;  #10 
a = 8'd209; b = 8'd90;  #10 
a = 8'd209; b = 8'd91;  #10 
a = 8'd209; b = 8'd92;  #10 
a = 8'd209; b = 8'd93;  #10 
a = 8'd209; b = 8'd94;  #10 
a = 8'd209; b = 8'd95;  #10 
a = 8'd209; b = 8'd96;  #10 
a = 8'd209; b = 8'd97;  #10 
a = 8'd209; b = 8'd98;  #10 
a = 8'd209; b = 8'd99;  #10 
a = 8'd209; b = 8'd100;  #10 
a = 8'd209; b = 8'd101;  #10 
a = 8'd209; b = 8'd102;  #10 
a = 8'd209; b = 8'd103;  #10 
a = 8'd209; b = 8'd104;  #10 
a = 8'd209; b = 8'd105;  #10 
a = 8'd209; b = 8'd106;  #10 
a = 8'd209; b = 8'd107;  #10 
a = 8'd209; b = 8'd108;  #10 
a = 8'd209; b = 8'd109;  #10 
a = 8'd209; b = 8'd110;  #10 
a = 8'd209; b = 8'd111;  #10 
a = 8'd209; b = 8'd112;  #10 
a = 8'd209; b = 8'd113;  #10 
a = 8'd209; b = 8'd114;  #10 
a = 8'd209; b = 8'd115;  #10 
a = 8'd209; b = 8'd116;  #10 
a = 8'd209; b = 8'd117;  #10 
a = 8'd209; b = 8'd118;  #10 
a = 8'd209; b = 8'd119;  #10 
a = 8'd209; b = 8'd120;  #10 
a = 8'd209; b = 8'd121;  #10 
a = 8'd209; b = 8'd122;  #10 
a = 8'd209; b = 8'd123;  #10 
a = 8'd209; b = 8'd124;  #10 
a = 8'd209; b = 8'd125;  #10 
a = 8'd209; b = 8'd126;  #10 
a = 8'd209; b = 8'd127;  #10 
a = 8'd209; b = 8'd128;  #10 
a = 8'd209; b = 8'd129;  #10 
a = 8'd209; b = 8'd130;  #10 
a = 8'd209; b = 8'd131;  #10 
a = 8'd209; b = 8'd132;  #10 
a = 8'd209; b = 8'd133;  #10 
a = 8'd209; b = 8'd134;  #10 
a = 8'd209; b = 8'd135;  #10 
a = 8'd209; b = 8'd136;  #10 
a = 8'd209; b = 8'd137;  #10 
a = 8'd209; b = 8'd138;  #10 
a = 8'd209; b = 8'd139;  #10 
a = 8'd209; b = 8'd140;  #10 
a = 8'd209; b = 8'd141;  #10 
a = 8'd209; b = 8'd142;  #10 
a = 8'd209; b = 8'd143;  #10 
a = 8'd209; b = 8'd144;  #10 
a = 8'd209; b = 8'd145;  #10 
a = 8'd209; b = 8'd146;  #10 
a = 8'd209; b = 8'd147;  #10 
a = 8'd209; b = 8'd148;  #10 
a = 8'd209; b = 8'd149;  #10 
a = 8'd209; b = 8'd150;  #10 
a = 8'd209; b = 8'd151;  #10 
a = 8'd209; b = 8'd152;  #10 
a = 8'd209; b = 8'd153;  #10 
a = 8'd209; b = 8'd154;  #10 
a = 8'd209; b = 8'd155;  #10 
a = 8'd209; b = 8'd156;  #10 
a = 8'd209; b = 8'd157;  #10 
a = 8'd209; b = 8'd158;  #10 
a = 8'd209; b = 8'd159;  #10 
a = 8'd209; b = 8'd160;  #10 
a = 8'd209; b = 8'd161;  #10 
a = 8'd209; b = 8'd162;  #10 
a = 8'd209; b = 8'd163;  #10 
a = 8'd209; b = 8'd164;  #10 
a = 8'd209; b = 8'd165;  #10 
a = 8'd209; b = 8'd166;  #10 
a = 8'd209; b = 8'd167;  #10 
a = 8'd209; b = 8'd168;  #10 
a = 8'd209; b = 8'd169;  #10 
a = 8'd209; b = 8'd170;  #10 
a = 8'd209; b = 8'd171;  #10 
a = 8'd209; b = 8'd172;  #10 
a = 8'd209; b = 8'd173;  #10 
a = 8'd209; b = 8'd174;  #10 
a = 8'd209; b = 8'd175;  #10 
a = 8'd209; b = 8'd176;  #10 
a = 8'd209; b = 8'd177;  #10 
a = 8'd209; b = 8'd178;  #10 
a = 8'd209; b = 8'd179;  #10 
a = 8'd209; b = 8'd180;  #10 
a = 8'd209; b = 8'd181;  #10 
a = 8'd209; b = 8'd182;  #10 
a = 8'd209; b = 8'd183;  #10 
a = 8'd209; b = 8'd184;  #10 
a = 8'd209; b = 8'd185;  #10 
a = 8'd209; b = 8'd186;  #10 
a = 8'd209; b = 8'd187;  #10 
a = 8'd209; b = 8'd188;  #10 
a = 8'd209; b = 8'd189;  #10 
a = 8'd209; b = 8'd190;  #10 
a = 8'd209; b = 8'd191;  #10 
a = 8'd209; b = 8'd192;  #10 
a = 8'd209; b = 8'd193;  #10 
a = 8'd209; b = 8'd194;  #10 
a = 8'd209; b = 8'd195;  #10 
a = 8'd209; b = 8'd196;  #10 
a = 8'd209; b = 8'd197;  #10 
a = 8'd209; b = 8'd198;  #10 
a = 8'd209; b = 8'd199;  #10 
a = 8'd209; b = 8'd200;  #10 
a = 8'd209; b = 8'd201;  #10 
a = 8'd209; b = 8'd202;  #10 
a = 8'd209; b = 8'd203;  #10 
a = 8'd209; b = 8'd204;  #10 
a = 8'd209; b = 8'd205;  #10 
a = 8'd209; b = 8'd206;  #10 
a = 8'd209; b = 8'd207;  #10 
a = 8'd209; b = 8'd208;  #10 
a = 8'd209; b = 8'd209;  #10 
a = 8'd209; b = 8'd210;  #10 
a = 8'd209; b = 8'd211;  #10 
a = 8'd209; b = 8'd212;  #10 
a = 8'd209; b = 8'd213;  #10 
a = 8'd209; b = 8'd214;  #10 
a = 8'd209; b = 8'd215;  #10 
a = 8'd209; b = 8'd216;  #10 
a = 8'd209; b = 8'd217;  #10 
a = 8'd209; b = 8'd218;  #10 
a = 8'd209; b = 8'd219;  #10 
a = 8'd209; b = 8'd220;  #10 
a = 8'd209; b = 8'd221;  #10 
a = 8'd209; b = 8'd222;  #10 
a = 8'd209; b = 8'd223;  #10 
a = 8'd209; b = 8'd224;  #10 
a = 8'd209; b = 8'd225;  #10 
a = 8'd209; b = 8'd226;  #10 
a = 8'd209; b = 8'd227;  #10 
a = 8'd209; b = 8'd228;  #10 
a = 8'd209; b = 8'd229;  #10 
a = 8'd209; b = 8'd230;  #10 
a = 8'd209; b = 8'd231;  #10 
a = 8'd209; b = 8'd232;  #10 
a = 8'd209; b = 8'd233;  #10 
a = 8'd209; b = 8'd234;  #10 
a = 8'd209; b = 8'd235;  #10 
a = 8'd209; b = 8'd236;  #10 
a = 8'd209; b = 8'd237;  #10 
a = 8'd209; b = 8'd238;  #10 
a = 8'd209; b = 8'd239;  #10 
a = 8'd209; b = 8'd240;  #10 
a = 8'd209; b = 8'd241;  #10 
a = 8'd209; b = 8'd242;  #10 
a = 8'd209; b = 8'd243;  #10 
a = 8'd209; b = 8'd244;  #10 
a = 8'd209; b = 8'd245;  #10 
a = 8'd209; b = 8'd246;  #10 
a = 8'd209; b = 8'd247;  #10 
a = 8'd209; b = 8'd248;  #10 
a = 8'd209; b = 8'd249;  #10 
a = 8'd209; b = 8'd250;  #10 
a = 8'd209; b = 8'd251;  #10 
a = 8'd209; b = 8'd252;  #10 
a = 8'd209; b = 8'd253;  #10 
a = 8'd209; b = 8'd254;  #10 
a = 8'd209; b = 8'd255;  #10 
a = 8'd210; b = 8'd0;  #10 
a = 8'd210; b = 8'd1;  #10 
a = 8'd210; b = 8'd2;  #10 
a = 8'd210; b = 8'd3;  #10 
a = 8'd210; b = 8'd4;  #10 
a = 8'd210; b = 8'd5;  #10 
a = 8'd210; b = 8'd6;  #10 
a = 8'd210; b = 8'd7;  #10 
a = 8'd210; b = 8'd8;  #10 
a = 8'd210; b = 8'd9;  #10 
a = 8'd210; b = 8'd10;  #10 
a = 8'd210; b = 8'd11;  #10 
a = 8'd210; b = 8'd12;  #10 
a = 8'd210; b = 8'd13;  #10 
a = 8'd210; b = 8'd14;  #10 
a = 8'd210; b = 8'd15;  #10 
a = 8'd210; b = 8'd16;  #10 
a = 8'd210; b = 8'd17;  #10 
a = 8'd210; b = 8'd18;  #10 
a = 8'd210; b = 8'd19;  #10 
a = 8'd210; b = 8'd20;  #10 
a = 8'd210; b = 8'd21;  #10 
a = 8'd210; b = 8'd22;  #10 
a = 8'd210; b = 8'd23;  #10 
a = 8'd210; b = 8'd24;  #10 
a = 8'd210; b = 8'd25;  #10 
a = 8'd210; b = 8'd26;  #10 
a = 8'd210; b = 8'd27;  #10 
a = 8'd210; b = 8'd28;  #10 
a = 8'd210; b = 8'd29;  #10 
a = 8'd210; b = 8'd30;  #10 
a = 8'd210; b = 8'd31;  #10 
a = 8'd210; b = 8'd32;  #10 
a = 8'd210; b = 8'd33;  #10 
a = 8'd210; b = 8'd34;  #10 
a = 8'd210; b = 8'd35;  #10 
a = 8'd210; b = 8'd36;  #10 
a = 8'd210; b = 8'd37;  #10 
a = 8'd210; b = 8'd38;  #10 
a = 8'd210; b = 8'd39;  #10 
a = 8'd210; b = 8'd40;  #10 
a = 8'd210; b = 8'd41;  #10 
a = 8'd210; b = 8'd42;  #10 
a = 8'd210; b = 8'd43;  #10 
a = 8'd210; b = 8'd44;  #10 
a = 8'd210; b = 8'd45;  #10 
a = 8'd210; b = 8'd46;  #10 
a = 8'd210; b = 8'd47;  #10 
a = 8'd210; b = 8'd48;  #10 
a = 8'd210; b = 8'd49;  #10 
a = 8'd210; b = 8'd50;  #10 
a = 8'd210; b = 8'd51;  #10 
a = 8'd210; b = 8'd52;  #10 
a = 8'd210; b = 8'd53;  #10 
a = 8'd210; b = 8'd54;  #10 
a = 8'd210; b = 8'd55;  #10 
a = 8'd210; b = 8'd56;  #10 
a = 8'd210; b = 8'd57;  #10 
a = 8'd210; b = 8'd58;  #10 
a = 8'd210; b = 8'd59;  #10 
a = 8'd210; b = 8'd60;  #10 
a = 8'd210; b = 8'd61;  #10 
a = 8'd210; b = 8'd62;  #10 
a = 8'd210; b = 8'd63;  #10 
a = 8'd210; b = 8'd64;  #10 
a = 8'd210; b = 8'd65;  #10 
a = 8'd210; b = 8'd66;  #10 
a = 8'd210; b = 8'd67;  #10 
a = 8'd210; b = 8'd68;  #10 
a = 8'd210; b = 8'd69;  #10 
a = 8'd210; b = 8'd70;  #10 
a = 8'd210; b = 8'd71;  #10 
a = 8'd210; b = 8'd72;  #10 
a = 8'd210; b = 8'd73;  #10 
a = 8'd210; b = 8'd74;  #10 
a = 8'd210; b = 8'd75;  #10 
a = 8'd210; b = 8'd76;  #10 
a = 8'd210; b = 8'd77;  #10 
a = 8'd210; b = 8'd78;  #10 
a = 8'd210; b = 8'd79;  #10 
a = 8'd210; b = 8'd80;  #10 
a = 8'd210; b = 8'd81;  #10 
a = 8'd210; b = 8'd82;  #10 
a = 8'd210; b = 8'd83;  #10 
a = 8'd210; b = 8'd84;  #10 
a = 8'd210; b = 8'd85;  #10 
a = 8'd210; b = 8'd86;  #10 
a = 8'd210; b = 8'd87;  #10 
a = 8'd210; b = 8'd88;  #10 
a = 8'd210; b = 8'd89;  #10 
a = 8'd210; b = 8'd90;  #10 
a = 8'd210; b = 8'd91;  #10 
a = 8'd210; b = 8'd92;  #10 
a = 8'd210; b = 8'd93;  #10 
a = 8'd210; b = 8'd94;  #10 
a = 8'd210; b = 8'd95;  #10 
a = 8'd210; b = 8'd96;  #10 
a = 8'd210; b = 8'd97;  #10 
a = 8'd210; b = 8'd98;  #10 
a = 8'd210; b = 8'd99;  #10 
a = 8'd210; b = 8'd100;  #10 
a = 8'd210; b = 8'd101;  #10 
a = 8'd210; b = 8'd102;  #10 
a = 8'd210; b = 8'd103;  #10 
a = 8'd210; b = 8'd104;  #10 
a = 8'd210; b = 8'd105;  #10 
a = 8'd210; b = 8'd106;  #10 
a = 8'd210; b = 8'd107;  #10 
a = 8'd210; b = 8'd108;  #10 
a = 8'd210; b = 8'd109;  #10 
a = 8'd210; b = 8'd110;  #10 
a = 8'd210; b = 8'd111;  #10 
a = 8'd210; b = 8'd112;  #10 
a = 8'd210; b = 8'd113;  #10 
a = 8'd210; b = 8'd114;  #10 
a = 8'd210; b = 8'd115;  #10 
a = 8'd210; b = 8'd116;  #10 
a = 8'd210; b = 8'd117;  #10 
a = 8'd210; b = 8'd118;  #10 
a = 8'd210; b = 8'd119;  #10 
a = 8'd210; b = 8'd120;  #10 
a = 8'd210; b = 8'd121;  #10 
a = 8'd210; b = 8'd122;  #10 
a = 8'd210; b = 8'd123;  #10 
a = 8'd210; b = 8'd124;  #10 
a = 8'd210; b = 8'd125;  #10 
a = 8'd210; b = 8'd126;  #10 
a = 8'd210; b = 8'd127;  #10 
a = 8'd210; b = 8'd128;  #10 
a = 8'd210; b = 8'd129;  #10 
a = 8'd210; b = 8'd130;  #10 
a = 8'd210; b = 8'd131;  #10 
a = 8'd210; b = 8'd132;  #10 
a = 8'd210; b = 8'd133;  #10 
a = 8'd210; b = 8'd134;  #10 
a = 8'd210; b = 8'd135;  #10 
a = 8'd210; b = 8'd136;  #10 
a = 8'd210; b = 8'd137;  #10 
a = 8'd210; b = 8'd138;  #10 
a = 8'd210; b = 8'd139;  #10 
a = 8'd210; b = 8'd140;  #10 
a = 8'd210; b = 8'd141;  #10 
a = 8'd210; b = 8'd142;  #10 
a = 8'd210; b = 8'd143;  #10 
a = 8'd210; b = 8'd144;  #10 
a = 8'd210; b = 8'd145;  #10 
a = 8'd210; b = 8'd146;  #10 
a = 8'd210; b = 8'd147;  #10 
a = 8'd210; b = 8'd148;  #10 
a = 8'd210; b = 8'd149;  #10 
a = 8'd210; b = 8'd150;  #10 
a = 8'd210; b = 8'd151;  #10 
a = 8'd210; b = 8'd152;  #10 
a = 8'd210; b = 8'd153;  #10 
a = 8'd210; b = 8'd154;  #10 
a = 8'd210; b = 8'd155;  #10 
a = 8'd210; b = 8'd156;  #10 
a = 8'd210; b = 8'd157;  #10 
a = 8'd210; b = 8'd158;  #10 
a = 8'd210; b = 8'd159;  #10 
a = 8'd210; b = 8'd160;  #10 
a = 8'd210; b = 8'd161;  #10 
a = 8'd210; b = 8'd162;  #10 
a = 8'd210; b = 8'd163;  #10 
a = 8'd210; b = 8'd164;  #10 
a = 8'd210; b = 8'd165;  #10 
a = 8'd210; b = 8'd166;  #10 
a = 8'd210; b = 8'd167;  #10 
a = 8'd210; b = 8'd168;  #10 
a = 8'd210; b = 8'd169;  #10 
a = 8'd210; b = 8'd170;  #10 
a = 8'd210; b = 8'd171;  #10 
a = 8'd210; b = 8'd172;  #10 
a = 8'd210; b = 8'd173;  #10 
a = 8'd210; b = 8'd174;  #10 
a = 8'd210; b = 8'd175;  #10 
a = 8'd210; b = 8'd176;  #10 
a = 8'd210; b = 8'd177;  #10 
a = 8'd210; b = 8'd178;  #10 
a = 8'd210; b = 8'd179;  #10 
a = 8'd210; b = 8'd180;  #10 
a = 8'd210; b = 8'd181;  #10 
a = 8'd210; b = 8'd182;  #10 
a = 8'd210; b = 8'd183;  #10 
a = 8'd210; b = 8'd184;  #10 
a = 8'd210; b = 8'd185;  #10 
a = 8'd210; b = 8'd186;  #10 
a = 8'd210; b = 8'd187;  #10 
a = 8'd210; b = 8'd188;  #10 
a = 8'd210; b = 8'd189;  #10 
a = 8'd210; b = 8'd190;  #10 
a = 8'd210; b = 8'd191;  #10 
a = 8'd210; b = 8'd192;  #10 
a = 8'd210; b = 8'd193;  #10 
a = 8'd210; b = 8'd194;  #10 
a = 8'd210; b = 8'd195;  #10 
a = 8'd210; b = 8'd196;  #10 
a = 8'd210; b = 8'd197;  #10 
a = 8'd210; b = 8'd198;  #10 
a = 8'd210; b = 8'd199;  #10 
a = 8'd210; b = 8'd200;  #10 
a = 8'd210; b = 8'd201;  #10 
a = 8'd210; b = 8'd202;  #10 
a = 8'd210; b = 8'd203;  #10 
a = 8'd210; b = 8'd204;  #10 
a = 8'd210; b = 8'd205;  #10 
a = 8'd210; b = 8'd206;  #10 
a = 8'd210; b = 8'd207;  #10 
a = 8'd210; b = 8'd208;  #10 
a = 8'd210; b = 8'd209;  #10 
a = 8'd210; b = 8'd210;  #10 
a = 8'd210; b = 8'd211;  #10 
a = 8'd210; b = 8'd212;  #10 
a = 8'd210; b = 8'd213;  #10 
a = 8'd210; b = 8'd214;  #10 
a = 8'd210; b = 8'd215;  #10 
a = 8'd210; b = 8'd216;  #10 
a = 8'd210; b = 8'd217;  #10 
a = 8'd210; b = 8'd218;  #10 
a = 8'd210; b = 8'd219;  #10 
a = 8'd210; b = 8'd220;  #10 
a = 8'd210; b = 8'd221;  #10 
a = 8'd210; b = 8'd222;  #10 
a = 8'd210; b = 8'd223;  #10 
a = 8'd210; b = 8'd224;  #10 
a = 8'd210; b = 8'd225;  #10 
a = 8'd210; b = 8'd226;  #10 
a = 8'd210; b = 8'd227;  #10 
a = 8'd210; b = 8'd228;  #10 
a = 8'd210; b = 8'd229;  #10 
a = 8'd210; b = 8'd230;  #10 
a = 8'd210; b = 8'd231;  #10 
a = 8'd210; b = 8'd232;  #10 
a = 8'd210; b = 8'd233;  #10 
a = 8'd210; b = 8'd234;  #10 
a = 8'd210; b = 8'd235;  #10 
a = 8'd210; b = 8'd236;  #10 
a = 8'd210; b = 8'd237;  #10 
a = 8'd210; b = 8'd238;  #10 
a = 8'd210; b = 8'd239;  #10 
a = 8'd210; b = 8'd240;  #10 
a = 8'd210; b = 8'd241;  #10 
a = 8'd210; b = 8'd242;  #10 
a = 8'd210; b = 8'd243;  #10 
a = 8'd210; b = 8'd244;  #10 
a = 8'd210; b = 8'd245;  #10 
a = 8'd210; b = 8'd246;  #10 
a = 8'd210; b = 8'd247;  #10 
a = 8'd210; b = 8'd248;  #10 
a = 8'd210; b = 8'd249;  #10 
a = 8'd210; b = 8'd250;  #10 
a = 8'd210; b = 8'd251;  #10 
a = 8'd210; b = 8'd252;  #10 
a = 8'd210; b = 8'd253;  #10 
a = 8'd210; b = 8'd254;  #10 
a = 8'd210; b = 8'd255;  #10 
a = 8'd211; b = 8'd0;  #10 
a = 8'd211; b = 8'd1;  #10 
a = 8'd211; b = 8'd2;  #10 
a = 8'd211; b = 8'd3;  #10 
a = 8'd211; b = 8'd4;  #10 
a = 8'd211; b = 8'd5;  #10 
a = 8'd211; b = 8'd6;  #10 
a = 8'd211; b = 8'd7;  #10 
a = 8'd211; b = 8'd8;  #10 
a = 8'd211; b = 8'd9;  #10 
a = 8'd211; b = 8'd10;  #10 
a = 8'd211; b = 8'd11;  #10 
a = 8'd211; b = 8'd12;  #10 
a = 8'd211; b = 8'd13;  #10 
a = 8'd211; b = 8'd14;  #10 
a = 8'd211; b = 8'd15;  #10 
a = 8'd211; b = 8'd16;  #10 
a = 8'd211; b = 8'd17;  #10 
a = 8'd211; b = 8'd18;  #10 
a = 8'd211; b = 8'd19;  #10 
a = 8'd211; b = 8'd20;  #10 
a = 8'd211; b = 8'd21;  #10 
a = 8'd211; b = 8'd22;  #10 
a = 8'd211; b = 8'd23;  #10 
a = 8'd211; b = 8'd24;  #10 
a = 8'd211; b = 8'd25;  #10 
a = 8'd211; b = 8'd26;  #10 
a = 8'd211; b = 8'd27;  #10 
a = 8'd211; b = 8'd28;  #10 
a = 8'd211; b = 8'd29;  #10 
a = 8'd211; b = 8'd30;  #10 
a = 8'd211; b = 8'd31;  #10 
a = 8'd211; b = 8'd32;  #10 
a = 8'd211; b = 8'd33;  #10 
a = 8'd211; b = 8'd34;  #10 
a = 8'd211; b = 8'd35;  #10 
a = 8'd211; b = 8'd36;  #10 
a = 8'd211; b = 8'd37;  #10 
a = 8'd211; b = 8'd38;  #10 
a = 8'd211; b = 8'd39;  #10 
a = 8'd211; b = 8'd40;  #10 
a = 8'd211; b = 8'd41;  #10 
a = 8'd211; b = 8'd42;  #10 
a = 8'd211; b = 8'd43;  #10 
a = 8'd211; b = 8'd44;  #10 
a = 8'd211; b = 8'd45;  #10 
a = 8'd211; b = 8'd46;  #10 
a = 8'd211; b = 8'd47;  #10 
a = 8'd211; b = 8'd48;  #10 
a = 8'd211; b = 8'd49;  #10 
a = 8'd211; b = 8'd50;  #10 
a = 8'd211; b = 8'd51;  #10 
a = 8'd211; b = 8'd52;  #10 
a = 8'd211; b = 8'd53;  #10 
a = 8'd211; b = 8'd54;  #10 
a = 8'd211; b = 8'd55;  #10 
a = 8'd211; b = 8'd56;  #10 
a = 8'd211; b = 8'd57;  #10 
a = 8'd211; b = 8'd58;  #10 
a = 8'd211; b = 8'd59;  #10 
a = 8'd211; b = 8'd60;  #10 
a = 8'd211; b = 8'd61;  #10 
a = 8'd211; b = 8'd62;  #10 
a = 8'd211; b = 8'd63;  #10 
a = 8'd211; b = 8'd64;  #10 
a = 8'd211; b = 8'd65;  #10 
a = 8'd211; b = 8'd66;  #10 
a = 8'd211; b = 8'd67;  #10 
a = 8'd211; b = 8'd68;  #10 
a = 8'd211; b = 8'd69;  #10 
a = 8'd211; b = 8'd70;  #10 
a = 8'd211; b = 8'd71;  #10 
a = 8'd211; b = 8'd72;  #10 
a = 8'd211; b = 8'd73;  #10 
a = 8'd211; b = 8'd74;  #10 
a = 8'd211; b = 8'd75;  #10 
a = 8'd211; b = 8'd76;  #10 
a = 8'd211; b = 8'd77;  #10 
a = 8'd211; b = 8'd78;  #10 
a = 8'd211; b = 8'd79;  #10 
a = 8'd211; b = 8'd80;  #10 
a = 8'd211; b = 8'd81;  #10 
a = 8'd211; b = 8'd82;  #10 
a = 8'd211; b = 8'd83;  #10 
a = 8'd211; b = 8'd84;  #10 
a = 8'd211; b = 8'd85;  #10 
a = 8'd211; b = 8'd86;  #10 
a = 8'd211; b = 8'd87;  #10 
a = 8'd211; b = 8'd88;  #10 
a = 8'd211; b = 8'd89;  #10 
a = 8'd211; b = 8'd90;  #10 
a = 8'd211; b = 8'd91;  #10 
a = 8'd211; b = 8'd92;  #10 
a = 8'd211; b = 8'd93;  #10 
a = 8'd211; b = 8'd94;  #10 
a = 8'd211; b = 8'd95;  #10 
a = 8'd211; b = 8'd96;  #10 
a = 8'd211; b = 8'd97;  #10 
a = 8'd211; b = 8'd98;  #10 
a = 8'd211; b = 8'd99;  #10 
a = 8'd211; b = 8'd100;  #10 
a = 8'd211; b = 8'd101;  #10 
a = 8'd211; b = 8'd102;  #10 
a = 8'd211; b = 8'd103;  #10 
a = 8'd211; b = 8'd104;  #10 
a = 8'd211; b = 8'd105;  #10 
a = 8'd211; b = 8'd106;  #10 
a = 8'd211; b = 8'd107;  #10 
a = 8'd211; b = 8'd108;  #10 
a = 8'd211; b = 8'd109;  #10 
a = 8'd211; b = 8'd110;  #10 
a = 8'd211; b = 8'd111;  #10 
a = 8'd211; b = 8'd112;  #10 
a = 8'd211; b = 8'd113;  #10 
a = 8'd211; b = 8'd114;  #10 
a = 8'd211; b = 8'd115;  #10 
a = 8'd211; b = 8'd116;  #10 
a = 8'd211; b = 8'd117;  #10 
a = 8'd211; b = 8'd118;  #10 
a = 8'd211; b = 8'd119;  #10 
a = 8'd211; b = 8'd120;  #10 
a = 8'd211; b = 8'd121;  #10 
a = 8'd211; b = 8'd122;  #10 
a = 8'd211; b = 8'd123;  #10 
a = 8'd211; b = 8'd124;  #10 
a = 8'd211; b = 8'd125;  #10 
a = 8'd211; b = 8'd126;  #10 
a = 8'd211; b = 8'd127;  #10 
a = 8'd211; b = 8'd128;  #10 
a = 8'd211; b = 8'd129;  #10 
a = 8'd211; b = 8'd130;  #10 
a = 8'd211; b = 8'd131;  #10 
a = 8'd211; b = 8'd132;  #10 
a = 8'd211; b = 8'd133;  #10 
a = 8'd211; b = 8'd134;  #10 
a = 8'd211; b = 8'd135;  #10 
a = 8'd211; b = 8'd136;  #10 
a = 8'd211; b = 8'd137;  #10 
a = 8'd211; b = 8'd138;  #10 
a = 8'd211; b = 8'd139;  #10 
a = 8'd211; b = 8'd140;  #10 
a = 8'd211; b = 8'd141;  #10 
a = 8'd211; b = 8'd142;  #10 
a = 8'd211; b = 8'd143;  #10 
a = 8'd211; b = 8'd144;  #10 
a = 8'd211; b = 8'd145;  #10 
a = 8'd211; b = 8'd146;  #10 
a = 8'd211; b = 8'd147;  #10 
a = 8'd211; b = 8'd148;  #10 
a = 8'd211; b = 8'd149;  #10 
a = 8'd211; b = 8'd150;  #10 
a = 8'd211; b = 8'd151;  #10 
a = 8'd211; b = 8'd152;  #10 
a = 8'd211; b = 8'd153;  #10 
a = 8'd211; b = 8'd154;  #10 
a = 8'd211; b = 8'd155;  #10 
a = 8'd211; b = 8'd156;  #10 
a = 8'd211; b = 8'd157;  #10 
a = 8'd211; b = 8'd158;  #10 
a = 8'd211; b = 8'd159;  #10 
a = 8'd211; b = 8'd160;  #10 
a = 8'd211; b = 8'd161;  #10 
a = 8'd211; b = 8'd162;  #10 
a = 8'd211; b = 8'd163;  #10 
a = 8'd211; b = 8'd164;  #10 
a = 8'd211; b = 8'd165;  #10 
a = 8'd211; b = 8'd166;  #10 
a = 8'd211; b = 8'd167;  #10 
a = 8'd211; b = 8'd168;  #10 
a = 8'd211; b = 8'd169;  #10 
a = 8'd211; b = 8'd170;  #10 
a = 8'd211; b = 8'd171;  #10 
a = 8'd211; b = 8'd172;  #10 
a = 8'd211; b = 8'd173;  #10 
a = 8'd211; b = 8'd174;  #10 
a = 8'd211; b = 8'd175;  #10 
a = 8'd211; b = 8'd176;  #10 
a = 8'd211; b = 8'd177;  #10 
a = 8'd211; b = 8'd178;  #10 
a = 8'd211; b = 8'd179;  #10 
a = 8'd211; b = 8'd180;  #10 
a = 8'd211; b = 8'd181;  #10 
a = 8'd211; b = 8'd182;  #10 
a = 8'd211; b = 8'd183;  #10 
a = 8'd211; b = 8'd184;  #10 
a = 8'd211; b = 8'd185;  #10 
a = 8'd211; b = 8'd186;  #10 
a = 8'd211; b = 8'd187;  #10 
a = 8'd211; b = 8'd188;  #10 
a = 8'd211; b = 8'd189;  #10 
a = 8'd211; b = 8'd190;  #10 
a = 8'd211; b = 8'd191;  #10 
a = 8'd211; b = 8'd192;  #10 
a = 8'd211; b = 8'd193;  #10 
a = 8'd211; b = 8'd194;  #10 
a = 8'd211; b = 8'd195;  #10 
a = 8'd211; b = 8'd196;  #10 
a = 8'd211; b = 8'd197;  #10 
a = 8'd211; b = 8'd198;  #10 
a = 8'd211; b = 8'd199;  #10 
a = 8'd211; b = 8'd200;  #10 
a = 8'd211; b = 8'd201;  #10 
a = 8'd211; b = 8'd202;  #10 
a = 8'd211; b = 8'd203;  #10 
a = 8'd211; b = 8'd204;  #10 
a = 8'd211; b = 8'd205;  #10 
a = 8'd211; b = 8'd206;  #10 
a = 8'd211; b = 8'd207;  #10 
a = 8'd211; b = 8'd208;  #10 
a = 8'd211; b = 8'd209;  #10 
a = 8'd211; b = 8'd210;  #10 
a = 8'd211; b = 8'd211;  #10 
a = 8'd211; b = 8'd212;  #10 
a = 8'd211; b = 8'd213;  #10 
a = 8'd211; b = 8'd214;  #10 
a = 8'd211; b = 8'd215;  #10 
a = 8'd211; b = 8'd216;  #10 
a = 8'd211; b = 8'd217;  #10 
a = 8'd211; b = 8'd218;  #10 
a = 8'd211; b = 8'd219;  #10 
a = 8'd211; b = 8'd220;  #10 
a = 8'd211; b = 8'd221;  #10 
a = 8'd211; b = 8'd222;  #10 
a = 8'd211; b = 8'd223;  #10 
a = 8'd211; b = 8'd224;  #10 
a = 8'd211; b = 8'd225;  #10 
a = 8'd211; b = 8'd226;  #10 
a = 8'd211; b = 8'd227;  #10 
a = 8'd211; b = 8'd228;  #10 
a = 8'd211; b = 8'd229;  #10 
a = 8'd211; b = 8'd230;  #10 
a = 8'd211; b = 8'd231;  #10 
a = 8'd211; b = 8'd232;  #10 
a = 8'd211; b = 8'd233;  #10 
a = 8'd211; b = 8'd234;  #10 
a = 8'd211; b = 8'd235;  #10 
a = 8'd211; b = 8'd236;  #10 
a = 8'd211; b = 8'd237;  #10 
a = 8'd211; b = 8'd238;  #10 
a = 8'd211; b = 8'd239;  #10 
a = 8'd211; b = 8'd240;  #10 
a = 8'd211; b = 8'd241;  #10 
a = 8'd211; b = 8'd242;  #10 
a = 8'd211; b = 8'd243;  #10 
a = 8'd211; b = 8'd244;  #10 
a = 8'd211; b = 8'd245;  #10 
a = 8'd211; b = 8'd246;  #10 
a = 8'd211; b = 8'd247;  #10 
a = 8'd211; b = 8'd248;  #10 
a = 8'd211; b = 8'd249;  #10 
a = 8'd211; b = 8'd250;  #10 
a = 8'd211; b = 8'd251;  #10 
a = 8'd211; b = 8'd252;  #10 
a = 8'd211; b = 8'd253;  #10 
a = 8'd211; b = 8'd254;  #10 
a = 8'd211; b = 8'd255;  #10 
a = 8'd212; b = 8'd0;  #10 
a = 8'd212; b = 8'd1;  #10 
a = 8'd212; b = 8'd2;  #10 
a = 8'd212; b = 8'd3;  #10 
a = 8'd212; b = 8'd4;  #10 
a = 8'd212; b = 8'd5;  #10 
a = 8'd212; b = 8'd6;  #10 
a = 8'd212; b = 8'd7;  #10 
a = 8'd212; b = 8'd8;  #10 
a = 8'd212; b = 8'd9;  #10 
a = 8'd212; b = 8'd10;  #10 
a = 8'd212; b = 8'd11;  #10 
a = 8'd212; b = 8'd12;  #10 
a = 8'd212; b = 8'd13;  #10 
a = 8'd212; b = 8'd14;  #10 
a = 8'd212; b = 8'd15;  #10 
a = 8'd212; b = 8'd16;  #10 
a = 8'd212; b = 8'd17;  #10 
a = 8'd212; b = 8'd18;  #10 
a = 8'd212; b = 8'd19;  #10 
a = 8'd212; b = 8'd20;  #10 
a = 8'd212; b = 8'd21;  #10 
a = 8'd212; b = 8'd22;  #10 
a = 8'd212; b = 8'd23;  #10 
a = 8'd212; b = 8'd24;  #10 
a = 8'd212; b = 8'd25;  #10 
a = 8'd212; b = 8'd26;  #10 
a = 8'd212; b = 8'd27;  #10 
a = 8'd212; b = 8'd28;  #10 
a = 8'd212; b = 8'd29;  #10 
a = 8'd212; b = 8'd30;  #10 
a = 8'd212; b = 8'd31;  #10 
a = 8'd212; b = 8'd32;  #10 
a = 8'd212; b = 8'd33;  #10 
a = 8'd212; b = 8'd34;  #10 
a = 8'd212; b = 8'd35;  #10 
a = 8'd212; b = 8'd36;  #10 
a = 8'd212; b = 8'd37;  #10 
a = 8'd212; b = 8'd38;  #10 
a = 8'd212; b = 8'd39;  #10 
a = 8'd212; b = 8'd40;  #10 
a = 8'd212; b = 8'd41;  #10 
a = 8'd212; b = 8'd42;  #10 
a = 8'd212; b = 8'd43;  #10 
a = 8'd212; b = 8'd44;  #10 
a = 8'd212; b = 8'd45;  #10 
a = 8'd212; b = 8'd46;  #10 
a = 8'd212; b = 8'd47;  #10 
a = 8'd212; b = 8'd48;  #10 
a = 8'd212; b = 8'd49;  #10 
a = 8'd212; b = 8'd50;  #10 
a = 8'd212; b = 8'd51;  #10 
a = 8'd212; b = 8'd52;  #10 
a = 8'd212; b = 8'd53;  #10 
a = 8'd212; b = 8'd54;  #10 
a = 8'd212; b = 8'd55;  #10 
a = 8'd212; b = 8'd56;  #10 
a = 8'd212; b = 8'd57;  #10 
a = 8'd212; b = 8'd58;  #10 
a = 8'd212; b = 8'd59;  #10 
a = 8'd212; b = 8'd60;  #10 
a = 8'd212; b = 8'd61;  #10 
a = 8'd212; b = 8'd62;  #10 
a = 8'd212; b = 8'd63;  #10 
a = 8'd212; b = 8'd64;  #10 
a = 8'd212; b = 8'd65;  #10 
a = 8'd212; b = 8'd66;  #10 
a = 8'd212; b = 8'd67;  #10 
a = 8'd212; b = 8'd68;  #10 
a = 8'd212; b = 8'd69;  #10 
a = 8'd212; b = 8'd70;  #10 
a = 8'd212; b = 8'd71;  #10 
a = 8'd212; b = 8'd72;  #10 
a = 8'd212; b = 8'd73;  #10 
a = 8'd212; b = 8'd74;  #10 
a = 8'd212; b = 8'd75;  #10 
a = 8'd212; b = 8'd76;  #10 
a = 8'd212; b = 8'd77;  #10 
a = 8'd212; b = 8'd78;  #10 
a = 8'd212; b = 8'd79;  #10 
a = 8'd212; b = 8'd80;  #10 
a = 8'd212; b = 8'd81;  #10 
a = 8'd212; b = 8'd82;  #10 
a = 8'd212; b = 8'd83;  #10 
a = 8'd212; b = 8'd84;  #10 
a = 8'd212; b = 8'd85;  #10 
a = 8'd212; b = 8'd86;  #10 
a = 8'd212; b = 8'd87;  #10 
a = 8'd212; b = 8'd88;  #10 
a = 8'd212; b = 8'd89;  #10 
a = 8'd212; b = 8'd90;  #10 
a = 8'd212; b = 8'd91;  #10 
a = 8'd212; b = 8'd92;  #10 
a = 8'd212; b = 8'd93;  #10 
a = 8'd212; b = 8'd94;  #10 
a = 8'd212; b = 8'd95;  #10 
a = 8'd212; b = 8'd96;  #10 
a = 8'd212; b = 8'd97;  #10 
a = 8'd212; b = 8'd98;  #10 
a = 8'd212; b = 8'd99;  #10 
a = 8'd212; b = 8'd100;  #10 
a = 8'd212; b = 8'd101;  #10 
a = 8'd212; b = 8'd102;  #10 
a = 8'd212; b = 8'd103;  #10 
a = 8'd212; b = 8'd104;  #10 
a = 8'd212; b = 8'd105;  #10 
a = 8'd212; b = 8'd106;  #10 
a = 8'd212; b = 8'd107;  #10 
a = 8'd212; b = 8'd108;  #10 
a = 8'd212; b = 8'd109;  #10 
a = 8'd212; b = 8'd110;  #10 
a = 8'd212; b = 8'd111;  #10 
a = 8'd212; b = 8'd112;  #10 
a = 8'd212; b = 8'd113;  #10 
a = 8'd212; b = 8'd114;  #10 
a = 8'd212; b = 8'd115;  #10 
a = 8'd212; b = 8'd116;  #10 
a = 8'd212; b = 8'd117;  #10 
a = 8'd212; b = 8'd118;  #10 
a = 8'd212; b = 8'd119;  #10 
a = 8'd212; b = 8'd120;  #10 
a = 8'd212; b = 8'd121;  #10 
a = 8'd212; b = 8'd122;  #10 
a = 8'd212; b = 8'd123;  #10 
a = 8'd212; b = 8'd124;  #10 
a = 8'd212; b = 8'd125;  #10 
a = 8'd212; b = 8'd126;  #10 
a = 8'd212; b = 8'd127;  #10 
a = 8'd212; b = 8'd128;  #10 
a = 8'd212; b = 8'd129;  #10 
a = 8'd212; b = 8'd130;  #10 
a = 8'd212; b = 8'd131;  #10 
a = 8'd212; b = 8'd132;  #10 
a = 8'd212; b = 8'd133;  #10 
a = 8'd212; b = 8'd134;  #10 
a = 8'd212; b = 8'd135;  #10 
a = 8'd212; b = 8'd136;  #10 
a = 8'd212; b = 8'd137;  #10 
a = 8'd212; b = 8'd138;  #10 
a = 8'd212; b = 8'd139;  #10 
a = 8'd212; b = 8'd140;  #10 
a = 8'd212; b = 8'd141;  #10 
a = 8'd212; b = 8'd142;  #10 
a = 8'd212; b = 8'd143;  #10 
a = 8'd212; b = 8'd144;  #10 
a = 8'd212; b = 8'd145;  #10 
a = 8'd212; b = 8'd146;  #10 
a = 8'd212; b = 8'd147;  #10 
a = 8'd212; b = 8'd148;  #10 
a = 8'd212; b = 8'd149;  #10 
a = 8'd212; b = 8'd150;  #10 
a = 8'd212; b = 8'd151;  #10 
a = 8'd212; b = 8'd152;  #10 
a = 8'd212; b = 8'd153;  #10 
a = 8'd212; b = 8'd154;  #10 
a = 8'd212; b = 8'd155;  #10 
a = 8'd212; b = 8'd156;  #10 
a = 8'd212; b = 8'd157;  #10 
a = 8'd212; b = 8'd158;  #10 
a = 8'd212; b = 8'd159;  #10 
a = 8'd212; b = 8'd160;  #10 
a = 8'd212; b = 8'd161;  #10 
a = 8'd212; b = 8'd162;  #10 
a = 8'd212; b = 8'd163;  #10 
a = 8'd212; b = 8'd164;  #10 
a = 8'd212; b = 8'd165;  #10 
a = 8'd212; b = 8'd166;  #10 
a = 8'd212; b = 8'd167;  #10 
a = 8'd212; b = 8'd168;  #10 
a = 8'd212; b = 8'd169;  #10 
a = 8'd212; b = 8'd170;  #10 
a = 8'd212; b = 8'd171;  #10 
a = 8'd212; b = 8'd172;  #10 
a = 8'd212; b = 8'd173;  #10 
a = 8'd212; b = 8'd174;  #10 
a = 8'd212; b = 8'd175;  #10 
a = 8'd212; b = 8'd176;  #10 
a = 8'd212; b = 8'd177;  #10 
a = 8'd212; b = 8'd178;  #10 
a = 8'd212; b = 8'd179;  #10 
a = 8'd212; b = 8'd180;  #10 
a = 8'd212; b = 8'd181;  #10 
a = 8'd212; b = 8'd182;  #10 
a = 8'd212; b = 8'd183;  #10 
a = 8'd212; b = 8'd184;  #10 
a = 8'd212; b = 8'd185;  #10 
a = 8'd212; b = 8'd186;  #10 
a = 8'd212; b = 8'd187;  #10 
a = 8'd212; b = 8'd188;  #10 
a = 8'd212; b = 8'd189;  #10 
a = 8'd212; b = 8'd190;  #10 
a = 8'd212; b = 8'd191;  #10 
a = 8'd212; b = 8'd192;  #10 
a = 8'd212; b = 8'd193;  #10 
a = 8'd212; b = 8'd194;  #10 
a = 8'd212; b = 8'd195;  #10 
a = 8'd212; b = 8'd196;  #10 
a = 8'd212; b = 8'd197;  #10 
a = 8'd212; b = 8'd198;  #10 
a = 8'd212; b = 8'd199;  #10 
a = 8'd212; b = 8'd200;  #10 
a = 8'd212; b = 8'd201;  #10 
a = 8'd212; b = 8'd202;  #10 
a = 8'd212; b = 8'd203;  #10 
a = 8'd212; b = 8'd204;  #10 
a = 8'd212; b = 8'd205;  #10 
a = 8'd212; b = 8'd206;  #10 
a = 8'd212; b = 8'd207;  #10 
a = 8'd212; b = 8'd208;  #10 
a = 8'd212; b = 8'd209;  #10 
a = 8'd212; b = 8'd210;  #10 
a = 8'd212; b = 8'd211;  #10 
a = 8'd212; b = 8'd212;  #10 
a = 8'd212; b = 8'd213;  #10 
a = 8'd212; b = 8'd214;  #10 
a = 8'd212; b = 8'd215;  #10 
a = 8'd212; b = 8'd216;  #10 
a = 8'd212; b = 8'd217;  #10 
a = 8'd212; b = 8'd218;  #10 
a = 8'd212; b = 8'd219;  #10 
a = 8'd212; b = 8'd220;  #10 
a = 8'd212; b = 8'd221;  #10 
a = 8'd212; b = 8'd222;  #10 
a = 8'd212; b = 8'd223;  #10 
a = 8'd212; b = 8'd224;  #10 
a = 8'd212; b = 8'd225;  #10 
a = 8'd212; b = 8'd226;  #10 
a = 8'd212; b = 8'd227;  #10 
a = 8'd212; b = 8'd228;  #10 
a = 8'd212; b = 8'd229;  #10 
a = 8'd212; b = 8'd230;  #10 
a = 8'd212; b = 8'd231;  #10 
a = 8'd212; b = 8'd232;  #10 
a = 8'd212; b = 8'd233;  #10 
a = 8'd212; b = 8'd234;  #10 
a = 8'd212; b = 8'd235;  #10 
a = 8'd212; b = 8'd236;  #10 
a = 8'd212; b = 8'd237;  #10 
a = 8'd212; b = 8'd238;  #10 
a = 8'd212; b = 8'd239;  #10 
a = 8'd212; b = 8'd240;  #10 
a = 8'd212; b = 8'd241;  #10 
a = 8'd212; b = 8'd242;  #10 
a = 8'd212; b = 8'd243;  #10 
a = 8'd212; b = 8'd244;  #10 
a = 8'd212; b = 8'd245;  #10 
a = 8'd212; b = 8'd246;  #10 
a = 8'd212; b = 8'd247;  #10 
a = 8'd212; b = 8'd248;  #10 
a = 8'd212; b = 8'd249;  #10 
a = 8'd212; b = 8'd250;  #10 
a = 8'd212; b = 8'd251;  #10 
a = 8'd212; b = 8'd252;  #10 
a = 8'd212; b = 8'd253;  #10 
a = 8'd212; b = 8'd254;  #10 
a = 8'd212; b = 8'd255;  #10 
a = 8'd213; b = 8'd0;  #10 
a = 8'd213; b = 8'd1;  #10 
a = 8'd213; b = 8'd2;  #10 
a = 8'd213; b = 8'd3;  #10 
a = 8'd213; b = 8'd4;  #10 
a = 8'd213; b = 8'd5;  #10 
a = 8'd213; b = 8'd6;  #10 
a = 8'd213; b = 8'd7;  #10 
a = 8'd213; b = 8'd8;  #10 
a = 8'd213; b = 8'd9;  #10 
a = 8'd213; b = 8'd10;  #10 
a = 8'd213; b = 8'd11;  #10 
a = 8'd213; b = 8'd12;  #10 
a = 8'd213; b = 8'd13;  #10 
a = 8'd213; b = 8'd14;  #10 
a = 8'd213; b = 8'd15;  #10 
a = 8'd213; b = 8'd16;  #10 
a = 8'd213; b = 8'd17;  #10 
a = 8'd213; b = 8'd18;  #10 
a = 8'd213; b = 8'd19;  #10 
a = 8'd213; b = 8'd20;  #10 
a = 8'd213; b = 8'd21;  #10 
a = 8'd213; b = 8'd22;  #10 
a = 8'd213; b = 8'd23;  #10 
a = 8'd213; b = 8'd24;  #10 
a = 8'd213; b = 8'd25;  #10 
a = 8'd213; b = 8'd26;  #10 
a = 8'd213; b = 8'd27;  #10 
a = 8'd213; b = 8'd28;  #10 
a = 8'd213; b = 8'd29;  #10 
a = 8'd213; b = 8'd30;  #10 
a = 8'd213; b = 8'd31;  #10 
a = 8'd213; b = 8'd32;  #10 
a = 8'd213; b = 8'd33;  #10 
a = 8'd213; b = 8'd34;  #10 
a = 8'd213; b = 8'd35;  #10 
a = 8'd213; b = 8'd36;  #10 
a = 8'd213; b = 8'd37;  #10 
a = 8'd213; b = 8'd38;  #10 
a = 8'd213; b = 8'd39;  #10 
a = 8'd213; b = 8'd40;  #10 
a = 8'd213; b = 8'd41;  #10 
a = 8'd213; b = 8'd42;  #10 
a = 8'd213; b = 8'd43;  #10 
a = 8'd213; b = 8'd44;  #10 
a = 8'd213; b = 8'd45;  #10 
a = 8'd213; b = 8'd46;  #10 
a = 8'd213; b = 8'd47;  #10 
a = 8'd213; b = 8'd48;  #10 
a = 8'd213; b = 8'd49;  #10 
a = 8'd213; b = 8'd50;  #10 
a = 8'd213; b = 8'd51;  #10 
a = 8'd213; b = 8'd52;  #10 
a = 8'd213; b = 8'd53;  #10 
a = 8'd213; b = 8'd54;  #10 
a = 8'd213; b = 8'd55;  #10 
a = 8'd213; b = 8'd56;  #10 
a = 8'd213; b = 8'd57;  #10 
a = 8'd213; b = 8'd58;  #10 
a = 8'd213; b = 8'd59;  #10 
a = 8'd213; b = 8'd60;  #10 
a = 8'd213; b = 8'd61;  #10 
a = 8'd213; b = 8'd62;  #10 
a = 8'd213; b = 8'd63;  #10 
a = 8'd213; b = 8'd64;  #10 
a = 8'd213; b = 8'd65;  #10 
a = 8'd213; b = 8'd66;  #10 
a = 8'd213; b = 8'd67;  #10 
a = 8'd213; b = 8'd68;  #10 
a = 8'd213; b = 8'd69;  #10 
a = 8'd213; b = 8'd70;  #10 
a = 8'd213; b = 8'd71;  #10 
a = 8'd213; b = 8'd72;  #10 
a = 8'd213; b = 8'd73;  #10 
a = 8'd213; b = 8'd74;  #10 
a = 8'd213; b = 8'd75;  #10 
a = 8'd213; b = 8'd76;  #10 
a = 8'd213; b = 8'd77;  #10 
a = 8'd213; b = 8'd78;  #10 
a = 8'd213; b = 8'd79;  #10 
a = 8'd213; b = 8'd80;  #10 
a = 8'd213; b = 8'd81;  #10 
a = 8'd213; b = 8'd82;  #10 
a = 8'd213; b = 8'd83;  #10 
a = 8'd213; b = 8'd84;  #10 
a = 8'd213; b = 8'd85;  #10 
a = 8'd213; b = 8'd86;  #10 
a = 8'd213; b = 8'd87;  #10 
a = 8'd213; b = 8'd88;  #10 
a = 8'd213; b = 8'd89;  #10 
a = 8'd213; b = 8'd90;  #10 
a = 8'd213; b = 8'd91;  #10 
a = 8'd213; b = 8'd92;  #10 
a = 8'd213; b = 8'd93;  #10 
a = 8'd213; b = 8'd94;  #10 
a = 8'd213; b = 8'd95;  #10 
a = 8'd213; b = 8'd96;  #10 
a = 8'd213; b = 8'd97;  #10 
a = 8'd213; b = 8'd98;  #10 
a = 8'd213; b = 8'd99;  #10 
a = 8'd213; b = 8'd100;  #10 
a = 8'd213; b = 8'd101;  #10 
a = 8'd213; b = 8'd102;  #10 
a = 8'd213; b = 8'd103;  #10 
a = 8'd213; b = 8'd104;  #10 
a = 8'd213; b = 8'd105;  #10 
a = 8'd213; b = 8'd106;  #10 
a = 8'd213; b = 8'd107;  #10 
a = 8'd213; b = 8'd108;  #10 
a = 8'd213; b = 8'd109;  #10 
a = 8'd213; b = 8'd110;  #10 
a = 8'd213; b = 8'd111;  #10 
a = 8'd213; b = 8'd112;  #10 
a = 8'd213; b = 8'd113;  #10 
a = 8'd213; b = 8'd114;  #10 
a = 8'd213; b = 8'd115;  #10 
a = 8'd213; b = 8'd116;  #10 
a = 8'd213; b = 8'd117;  #10 
a = 8'd213; b = 8'd118;  #10 
a = 8'd213; b = 8'd119;  #10 
a = 8'd213; b = 8'd120;  #10 
a = 8'd213; b = 8'd121;  #10 
a = 8'd213; b = 8'd122;  #10 
a = 8'd213; b = 8'd123;  #10 
a = 8'd213; b = 8'd124;  #10 
a = 8'd213; b = 8'd125;  #10 
a = 8'd213; b = 8'd126;  #10 
a = 8'd213; b = 8'd127;  #10 
a = 8'd213; b = 8'd128;  #10 
a = 8'd213; b = 8'd129;  #10 
a = 8'd213; b = 8'd130;  #10 
a = 8'd213; b = 8'd131;  #10 
a = 8'd213; b = 8'd132;  #10 
a = 8'd213; b = 8'd133;  #10 
a = 8'd213; b = 8'd134;  #10 
a = 8'd213; b = 8'd135;  #10 
a = 8'd213; b = 8'd136;  #10 
a = 8'd213; b = 8'd137;  #10 
a = 8'd213; b = 8'd138;  #10 
a = 8'd213; b = 8'd139;  #10 
a = 8'd213; b = 8'd140;  #10 
a = 8'd213; b = 8'd141;  #10 
a = 8'd213; b = 8'd142;  #10 
a = 8'd213; b = 8'd143;  #10 
a = 8'd213; b = 8'd144;  #10 
a = 8'd213; b = 8'd145;  #10 
a = 8'd213; b = 8'd146;  #10 
a = 8'd213; b = 8'd147;  #10 
a = 8'd213; b = 8'd148;  #10 
a = 8'd213; b = 8'd149;  #10 
a = 8'd213; b = 8'd150;  #10 
a = 8'd213; b = 8'd151;  #10 
a = 8'd213; b = 8'd152;  #10 
a = 8'd213; b = 8'd153;  #10 
a = 8'd213; b = 8'd154;  #10 
a = 8'd213; b = 8'd155;  #10 
a = 8'd213; b = 8'd156;  #10 
a = 8'd213; b = 8'd157;  #10 
a = 8'd213; b = 8'd158;  #10 
a = 8'd213; b = 8'd159;  #10 
a = 8'd213; b = 8'd160;  #10 
a = 8'd213; b = 8'd161;  #10 
a = 8'd213; b = 8'd162;  #10 
a = 8'd213; b = 8'd163;  #10 
a = 8'd213; b = 8'd164;  #10 
a = 8'd213; b = 8'd165;  #10 
a = 8'd213; b = 8'd166;  #10 
a = 8'd213; b = 8'd167;  #10 
a = 8'd213; b = 8'd168;  #10 
a = 8'd213; b = 8'd169;  #10 
a = 8'd213; b = 8'd170;  #10 
a = 8'd213; b = 8'd171;  #10 
a = 8'd213; b = 8'd172;  #10 
a = 8'd213; b = 8'd173;  #10 
a = 8'd213; b = 8'd174;  #10 
a = 8'd213; b = 8'd175;  #10 
a = 8'd213; b = 8'd176;  #10 
a = 8'd213; b = 8'd177;  #10 
a = 8'd213; b = 8'd178;  #10 
a = 8'd213; b = 8'd179;  #10 
a = 8'd213; b = 8'd180;  #10 
a = 8'd213; b = 8'd181;  #10 
a = 8'd213; b = 8'd182;  #10 
a = 8'd213; b = 8'd183;  #10 
a = 8'd213; b = 8'd184;  #10 
a = 8'd213; b = 8'd185;  #10 
a = 8'd213; b = 8'd186;  #10 
a = 8'd213; b = 8'd187;  #10 
a = 8'd213; b = 8'd188;  #10 
a = 8'd213; b = 8'd189;  #10 
a = 8'd213; b = 8'd190;  #10 
a = 8'd213; b = 8'd191;  #10 
a = 8'd213; b = 8'd192;  #10 
a = 8'd213; b = 8'd193;  #10 
a = 8'd213; b = 8'd194;  #10 
a = 8'd213; b = 8'd195;  #10 
a = 8'd213; b = 8'd196;  #10 
a = 8'd213; b = 8'd197;  #10 
a = 8'd213; b = 8'd198;  #10 
a = 8'd213; b = 8'd199;  #10 
a = 8'd213; b = 8'd200;  #10 
a = 8'd213; b = 8'd201;  #10 
a = 8'd213; b = 8'd202;  #10 
a = 8'd213; b = 8'd203;  #10 
a = 8'd213; b = 8'd204;  #10 
a = 8'd213; b = 8'd205;  #10 
a = 8'd213; b = 8'd206;  #10 
a = 8'd213; b = 8'd207;  #10 
a = 8'd213; b = 8'd208;  #10 
a = 8'd213; b = 8'd209;  #10 
a = 8'd213; b = 8'd210;  #10 
a = 8'd213; b = 8'd211;  #10 
a = 8'd213; b = 8'd212;  #10 
a = 8'd213; b = 8'd213;  #10 
a = 8'd213; b = 8'd214;  #10 
a = 8'd213; b = 8'd215;  #10 
a = 8'd213; b = 8'd216;  #10 
a = 8'd213; b = 8'd217;  #10 
a = 8'd213; b = 8'd218;  #10 
a = 8'd213; b = 8'd219;  #10 
a = 8'd213; b = 8'd220;  #10 
a = 8'd213; b = 8'd221;  #10 
a = 8'd213; b = 8'd222;  #10 
a = 8'd213; b = 8'd223;  #10 
a = 8'd213; b = 8'd224;  #10 
a = 8'd213; b = 8'd225;  #10 
a = 8'd213; b = 8'd226;  #10 
a = 8'd213; b = 8'd227;  #10 
a = 8'd213; b = 8'd228;  #10 
a = 8'd213; b = 8'd229;  #10 
a = 8'd213; b = 8'd230;  #10 
a = 8'd213; b = 8'd231;  #10 
a = 8'd213; b = 8'd232;  #10 
a = 8'd213; b = 8'd233;  #10 
a = 8'd213; b = 8'd234;  #10 
a = 8'd213; b = 8'd235;  #10 
a = 8'd213; b = 8'd236;  #10 
a = 8'd213; b = 8'd237;  #10 
a = 8'd213; b = 8'd238;  #10 
a = 8'd213; b = 8'd239;  #10 
a = 8'd213; b = 8'd240;  #10 
a = 8'd213; b = 8'd241;  #10 
a = 8'd213; b = 8'd242;  #10 
a = 8'd213; b = 8'd243;  #10 
a = 8'd213; b = 8'd244;  #10 
a = 8'd213; b = 8'd245;  #10 
a = 8'd213; b = 8'd246;  #10 
a = 8'd213; b = 8'd247;  #10 
a = 8'd213; b = 8'd248;  #10 
a = 8'd213; b = 8'd249;  #10 
a = 8'd213; b = 8'd250;  #10 
a = 8'd213; b = 8'd251;  #10 
a = 8'd213; b = 8'd252;  #10 
a = 8'd213; b = 8'd253;  #10 
a = 8'd213; b = 8'd254;  #10 
a = 8'd213; b = 8'd255;  #10 
a = 8'd214; b = 8'd0;  #10 
a = 8'd214; b = 8'd1;  #10 
a = 8'd214; b = 8'd2;  #10 
a = 8'd214; b = 8'd3;  #10 
a = 8'd214; b = 8'd4;  #10 
a = 8'd214; b = 8'd5;  #10 
a = 8'd214; b = 8'd6;  #10 
a = 8'd214; b = 8'd7;  #10 
a = 8'd214; b = 8'd8;  #10 
a = 8'd214; b = 8'd9;  #10 
a = 8'd214; b = 8'd10;  #10 
a = 8'd214; b = 8'd11;  #10 
a = 8'd214; b = 8'd12;  #10 
a = 8'd214; b = 8'd13;  #10 
a = 8'd214; b = 8'd14;  #10 
a = 8'd214; b = 8'd15;  #10 
a = 8'd214; b = 8'd16;  #10 
a = 8'd214; b = 8'd17;  #10 
a = 8'd214; b = 8'd18;  #10 
a = 8'd214; b = 8'd19;  #10 
a = 8'd214; b = 8'd20;  #10 
a = 8'd214; b = 8'd21;  #10 
a = 8'd214; b = 8'd22;  #10 
a = 8'd214; b = 8'd23;  #10 
a = 8'd214; b = 8'd24;  #10 
a = 8'd214; b = 8'd25;  #10 
a = 8'd214; b = 8'd26;  #10 
a = 8'd214; b = 8'd27;  #10 
a = 8'd214; b = 8'd28;  #10 
a = 8'd214; b = 8'd29;  #10 
a = 8'd214; b = 8'd30;  #10 
a = 8'd214; b = 8'd31;  #10 
a = 8'd214; b = 8'd32;  #10 
a = 8'd214; b = 8'd33;  #10 
a = 8'd214; b = 8'd34;  #10 
a = 8'd214; b = 8'd35;  #10 
a = 8'd214; b = 8'd36;  #10 
a = 8'd214; b = 8'd37;  #10 
a = 8'd214; b = 8'd38;  #10 
a = 8'd214; b = 8'd39;  #10 
a = 8'd214; b = 8'd40;  #10 
a = 8'd214; b = 8'd41;  #10 
a = 8'd214; b = 8'd42;  #10 
a = 8'd214; b = 8'd43;  #10 
a = 8'd214; b = 8'd44;  #10 
a = 8'd214; b = 8'd45;  #10 
a = 8'd214; b = 8'd46;  #10 
a = 8'd214; b = 8'd47;  #10 
a = 8'd214; b = 8'd48;  #10 
a = 8'd214; b = 8'd49;  #10 
a = 8'd214; b = 8'd50;  #10 
a = 8'd214; b = 8'd51;  #10 
a = 8'd214; b = 8'd52;  #10 
a = 8'd214; b = 8'd53;  #10 
a = 8'd214; b = 8'd54;  #10 
a = 8'd214; b = 8'd55;  #10 
a = 8'd214; b = 8'd56;  #10 
a = 8'd214; b = 8'd57;  #10 
a = 8'd214; b = 8'd58;  #10 
a = 8'd214; b = 8'd59;  #10 
a = 8'd214; b = 8'd60;  #10 
a = 8'd214; b = 8'd61;  #10 
a = 8'd214; b = 8'd62;  #10 
a = 8'd214; b = 8'd63;  #10 
a = 8'd214; b = 8'd64;  #10 
a = 8'd214; b = 8'd65;  #10 
a = 8'd214; b = 8'd66;  #10 
a = 8'd214; b = 8'd67;  #10 
a = 8'd214; b = 8'd68;  #10 
a = 8'd214; b = 8'd69;  #10 
a = 8'd214; b = 8'd70;  #10 
a = 8'd214; b = 8'd71;  #10 
a = 8'd214; b = 8'd72;  #10 
a = 8'd214; b = 8'd73;  #10 
a = 8'd214; b = 8'd74;  #10 
a = 8'd214; b = 8'd75;  #10 
a = 8'd214; b = 8'd76;  #10 
a = 8'd214; b = 8'd77;  #10 
a = 8'd214; b = 8'd78;  #10 
a = 8'd214; b = 8'd79;  #10 
a = 8'd214; b = 8'd80;  #10 
a = 8'd214; b = 8'd81;  #10 
a = 8'd214; b = 8'd82;  #10 
a = 8'd214; b = 8'd83;  #10 
a = 8'd214; b = 8'd84;  #10 
a = 8'd214; b = 8'd85;  #10 
a = 8'd214; b = 8'd86;  #10 
a = 8'd214; b = 8'd87;  #10 
a = 8'd214; b = 8'd88;  #10 
a = 8'd214; b = 8'd89;  #10 
a = 8'd214; b = 8'd90;  #10 
a = 8'd214; b = 8'd91;  #10 
a = 8'd214; b = 8'd92;  #10 
a = 8'd214; b = 8'd93;  #10 
a = 8'd214; b = 8'd94;  #10 
a = 8'd214; b = 8'd95;  #10 
a = 8'd214; b = 8'd96;  #10 
a = 8'd214; b = 8'd97;  #10 
a = 8'd214; b = 8'd98;  #10 
a = 8'd214; b = 8'd99;  #10 
a = 8'd214; b = 8'd100;  #10 
a = 8'd214; b = 8'd101;  #10 
a = 8'd214; b = 8'd102;  #10 
a = 8'd214; b = 8'd103;  #10 
a = 8'd214; b = 8'd104;  #10 
a = 8'd214; b = 8'd105;  #10 
a = 8'd214; b = 8'd106;  #10 
a = 8'd214; b = 8'd107;  #10 
a = 8'd214; b = 8'd108;  #10 
a = 8'd214; b = 8'd109;  #10 
a = 8'd214; b = 8'd110;  #10 
a = 8'd214; b = 8'd111;  #10 
a = 8'd214; b = 8'd112;  #10 
a = 8'd214; b = 8'd113;  #10 
a = 8'd214; b = 8'd114;  #10 
a = 8'd214; b = 8'd115;  #10 
a = 8'd214; b = 8'd116;  #10 
a = 8'd214; b = 8'd117;  #10 
a = 8'd214; b = 8'd118;  #10 
a = 8'd214; b = 8'd119;  #10 
a = 8'd214; b = 8'd120;  #10 
a = 8'd214; b = 8'd121;  #10 
a = 8'd214; b = 8'd122;  #10 
a = 8'd214; b = 8'd123;  #10 
a = 8'd214; b = 8'd124;  #10 
a = 8'd214; b = 8'd125;  #10 
a = 8'd214; b = 8'd126;  #10 
a = 8'd214; b = 8'd127;  #10 
a = 8'd214; b = 8'd128;  #10 
a = 8'd214; b = 8'd129;  #10 
a = 8'd214; b = 8'd130;  #10 
a = 8'd214; b = 8'd131;  #10 
a = 8'd214; b = 8'd132;  #10 
a = 8'd214; b = 8'd133;  #10 
a = 8'd214; b = 8'd134;  #10 
a = 8'd214; b = 8'd135;  #10 
a = 8'd214; b = 8'd136;  #10 
a = 8'd214; b = 8'd137;  #10 
a = 8'd214; b = 8'd138;  #10 
a = 8'd214; b = 8'd139;  #10 
a = 8'd214; b = 8'd140;  #10 
a = 8'd214; b = 8'd141;  #10 
a = 8'd214; b = 8'd142;  #10 
a = 8'd214; b = 8'd143;  #10 
a = 8'd214; b = 8'd144;  #10 
a = 8'd214; b = 8'd145;  #10 
a = 8'd214; b = 8'd146;  #10 
a = 8'd214; b = 8'd147;  #10 
a = 8'd214; b = 8'd148;  #10 
a = 8'd214; b = 8'd149;  #10 
a = 8'd214; b = 8'd150;  #10 
a = 8'd214; b = 8'd151;  #10 
a = 8'd214; b = 8'd152;  #10 
a = 8'd214; b = 8'd153;  #10 
a = 8'd214; b = 8'd154;  #10 
a = 8'd214; b = 8'd155;  #10 
a = 8'd214; b = 8'd156;  #10 
a = 8'd214; b = 8'd157;  #10 
a = 8'd214; b = 8'd158;  #10 
a = 8'd214; b = 8'd159;  #10 
a = 8'd214; b = 8'd160;  #10 
a = 8'd214; b = 8'd161;  #10 
a = 8'd214; b = 8'd162;  #10 
a = 8'd214; b = 8'd163;  #10 
a = 8'd214; b = 8'd164;  #10 
a = 8'd214; b = 8'd165;  #10 
a = 8'd214; b = 8'd166;  #10 
a = 8'd214; b = 8'd167;  #10 
a = 8'd214; b = 8'd168;  #10 
a = 8'd214; b = 8'd169;  #10 
a = 8'd214; b = 8'd170;  #10 
a = 8'd214; b = 8'd171;  #10 
a = 8'd214; b = 8'd172;  #10 
a = 8'd214; b = 8'd173;  #10 
a = 8'd214; b = 8'd174;  #10 
a = 8'd214; b = 8'd175;  #10 
a = 8'd214; b = 8'd176;  #10 
a = 8'd214; b = 8'd177;  #10 
a = 8'd214; b = 8'd178;  #10 
a = 8'd214; b = 8'd179;  #10 
a = 8'd214; b = 8'd180;  #10 
a = 8'd214; b = 8'd181;  #10 
a = 8'd214; b = 8'd182;  #10 
a = 8'd214; b = 8'd183;  #10 
a = 8'd214; b = 8'd184;  #10 
a = 8'd214; b = 8'd185;  #10 
a = 8'd214; b = 8'd186;  #10 
a = 8'd214; b = 8'd187;  #10 
a = 8'd214; b = 8'd188;  #10 
a = 8'd214; b = 8'd189;  #10 
a = 8'd214; b = 8'd190;  #10 
a = 8'd214; b = 8'd191;  #10 
a = 8'd214; b = 8'd192;  #10 
a = 8'd214; b = 8'd193;  #10 
a = 8'd214; b = 8'd194;  #10 
a = 8'd214; b = 8'd195;  #10 
a = 8'd214; b = 8'd196;  #10 
a = 8'd214; b = 8'd197;  #10 
a = 8'd214; b = 8'd198;  #10 
a = 8'd214; b = 8'd199;  #10 
a = 8'd214; b = 8'd200;  #10 
a = 8'd214; b = 8'd201;  #10 
a = 8'd214; b = 8'd202;  #10 
a = 8'd214; b = 8'd203;  #10 
a = 8'd214; b = 8'd204;  #10 
a = 8'd214; b = 8'd205;  #10 
a = 8'd214; b = 8'd206;  #10 
a = 8'd214; b = 8'd207;  #10 
a = 8'd214; b = 8'd208;  #10 
a = 8'd214; b = 8'd209;  #10 
a = 8'd214; b = 8'd210;  #10 
a = 8'd214; b = 8'd211;  #10 
a = 8'd214; b = 8'd212;  #10 
a = 8'd214; b = 8'd213;  #10 
a = 8'd214; b = 8'd214;  #10 
a = 8'd214; b = 8'd215;  #10 
a = 8'd214; b = 8'd216;  #10 
a = 8'd214; b = 8'd217;  #10 
a = 8'd214; b = 8'd218;  #10 
a = 8'd214; b = 8'd219;  #10 
a = 8'd214; b = 8'd220;  #10 
a = 8'd214; b = 8'd221;  #10 
a = 8'd214; b = 8'd222;  #10 
a = 8'd214; b = 8'd223;  #10 
a = 8'd214; b = 8'd224;  #10 
a = 8'd214; b = 8'd225;  #10 
a = 8'd214; b = 8'd226;  #10 
a = 8'd214; b = 8'd227;  #10 
a = 8'd214; b = 8'd228;  #10 
a = 8'd214; b = 8'd229;  #10 
a = 8'd214; b = 8'd230;  #10 
a = 8'd214; b = 8'd231;  #10 
a = 8'd214; b = 8'd232;  #10 
a = 8'd214; b = 8'd233;  #10 
a = 8'd214; b = 8'd234;  #10 
a = 8'd214; b = 8'd235;  #10 
a = 8'd214; b = 8'd236;  #10 
a = 8'd214; b = 8'd237;  #10 
a = 8'd214; b = 8'd238;  #10 
a = 8'd214; b = 8'd239;  #10 
a = 8'd214; b = 8'd240;  #10 
a = 8'd214; b = 8'd241;  #10 
a = 8'd214; b = 8'd242;  #10 
a = 8'd214; b = 8'd243;  #10 
a = 8'd214; b = 8'd244;  #10 
a = 8'd214; b = 8'd245;  #10 
a = 8'd214; b = 8'd246;  #10 
a = 8'd214; b = 8'd247;  #10 
a = 8'd214; b = 8'd248;  #10 
a = 8'd214; b = 8'd249;  #10 
a = 8'd214; b = 8'd250;  #10 
a = 8'd214; b = 8'd251;  #10 
a = 8'd214; b = 8'd252;  #10 
a = 8'd214; b = 8'd253;  #10 
a = 8'd214; b = 8'd254;  #10 
a = 8'd214; b = 8'd255;  #10 
a = 8'd215; b = 8'd0;  #10 
a = 8'd215; b = 8'd1;  #10 
a = 8'd215; b = 8'd2;  #10 
a = 8'd215; b = 8'd3;  #10 
a = 8'd215; b = 8'd4;  #10 
a = 8'd215; b = 8'd5;  #10 
a = 8'd215; b = 8'd6;  #10 
a = 8'd215; b = 8'd7;  #10 
a = 8'd215; b = 8'd8;  #10 
a = 8'd215; b = 8'd9;  #10 
a = 8'd215; b = 8'd10;  #10 
a = 8'd215; b = 8'd11;  #10 
a = 8'd215; b = 8'd12;  #10 
a = 8'd215; b = 8'd13;  #10 
a = 8'd215; b = 8'd14;  #10 
a = 8'd215; b = 8'd15;  #10 
a = 8'd215; b = 8'd16;  #10 
a = 8'd215; b = 8'd17;  #10 
a = 8'd215; b = 8'd18;  #10 
a = 8'd215; b = 8'd19;  #10 
a = 8'd215; b = 8'd20;  #10 
a = 8'd215; b = 8'd21;  #10 
a = 8'd215; b = 8'd22;  #10 
a = 8'd215; b = 8'd23;  #10 
a = 8'd215; b = 8'd24;  #10 
a = 8'd215; b = 8'd25;  #10 
a = 8'd215; b = 8'd26;  #10 
a = 8'd215; b = 8'd27;  #10 
a = 8'd215; b = 8'd28;  #10 
a = 8'd215; b = 8'd29;  #10 
a = 8'd215; b = 8'd30;  #10 
a = 8'd215; b = 8'd31;  #10 
a = 8'd215; b = 8'd32;  #10 
a = 8'd215; b = 8'd33;  #10 
a = 8'd215; b = 8'd34;  #10 
a = 8'd215; b = 8'd35;  #10 
a = 8'd215; b = 8'd36;  #10 
a = 8'd215; b = 8'd37;  #10 
a = 8'd215; b = 8'd38;  #10 
a = 8'd215; b = 8'd39;  #10 
a = 8'd215; b = 8'd40;  #10 
a = 8'd215; b = 8'd41;  #10 
a = 8'd215; b = 8'd42;  #10 
a = 8'd215; b = 8'd43;  #10 
a = 8'd215; b = 8'd44;  #10 
a = 8'd215; b = 8'd45;  #10 
a = 8'd215; b = 8'd46;  #10 
a = 8'd215; b = 8'd47;  #10 
a = 8'd215; b = 8'd48;  #10 
a = 8'd215; b = 8'd49;  #10 
a = 8'd215; b = 8'd50;  #10 
a = 8'd215; b = 8'd51;  #10 
a = 8'd215; b = 8'd52;  #10 
a = 8'd215; b = 8'd53;  #10 
a = 8'd215; b = 8'd54;  #10 
a = 8'd215; b = 8'd55;  #10 
a = 8'd215; b = 8'd56;  #10 
a = 8'd215; b = 8'd57;  #10 
a = 8'd215; b = 8'd58;  #10 
a = 8'd215; b = 8'd59;  #10 
a = 8'd215; b = 8'd60;  #10 
a = 8'd215; b = 8'd61;  #10 
a = 8'd215; b = 8'd62;  #10 
a = 8'd215; b = 8'd63;  #10 
a = 8'd215; b = 8'd64;  #10 
a = 8'd215; b = 8'd65;  #10 
a = 8'd215; b = 8'd66;  #10 
a = 8'd215; b = 8'd67;  #10 
a = 8'd215; b = 8'd68;  #10 
a = 8'd215; b = 8'd69;  #10 
a = 8'd215; b = 8'd70;  #10 
a = 8'd215; b = 8'd71;  #10 
a = 8'd215; b = 8'd72;  #10 
a = 8'd215; b = 8'd73;  #10 
a = 8'd215; b = 8'd74;  #10 
a = 8'd215; b = 8'd75;  #10 
a = 8'd215; b = 8'd76;  #10 
a = 8'd215; b = 8'd77;  #10 
a = 8'd215; b = 8'd78;  #10 
a = 8'd215; b = 8'd79;  #10 
a = 8'd215; b = 8'd80;  #10 
a = 8'd215; b = 8'd81;  #10 
a = 8'd215; b = 8'd82;  #10 
a = 8'd215; b = 8'd83;  #10 
a = 8'd215; b = 8'd84;  #10 
a = 8'd215; b = 8'd85;  #10 
a = 8'd215; b = 8'd86;  #10 
a = 8'd215; b = 8'd87;  #10 
a = 8'd215; b = 8'd88;  #10 
a = 8'd215; b = 8'd89;  #10 
a = 8'd215; b = 8'd90;  #10 
a = 8'd215; b = 8'd91;  #10 
a = 8'd215; b = 8'd92;  #10 
a = 8'd215; b = 8'd93;  #10 
a = 8'd215; b = 8'd94;  #10 
a = 8'd215; b = 8'd95;  #10 
a = 8'd215; b = 8'd96;  #10 
a = 8'd215; b = 8'd97;  #10 
a = 8'd215; b = 8'd98;  #10 
a = 8'd215; b = 8'd99;  #10 
a = 8'd215; b = 8'd100;  #10 
a = 8'd215; b = 8'd101;  #10 
a = 8'd215; b = 8'd102;  #10 
a = 8'd215; b = 8'd103;  #10 
a = 8'd215; b = 8'd104;  #10 
a = 8'd215; b = 8'd105;  #10 
a = 8'd215; b = 8'd106;  #10 
a = 8'd215; b = 8'd107;  #10 
a = 8'd215; b = 8'd108;  #10 
a = 8'd215; b = 8'd109;  #10 
a = 8'd215; b = 8'd110;  #10 
a = 8'd215; b = 8'd111;  #10 
a = 8'd215; b = 8'd112;  #10 
a = 8'd215; b = 8'd113;  #10 
a = 8'd215; b = 8'd114;  #10 
a = 8'd215; b = 8'd115;  #10 
a = 8'd215; b = 8'd116;  #10 
a = 8'd215; b = 8'd117;  #10 
a = 8'd215; b = 8'd118;  #10 
a = 8'd215; b = 8'd119;  #10 
a = 8'd215; b = 8'd120;  #10 
a = 8'd215; b = 8'd121;  #10 
a = 8'd215; b = 8'd122;  #10 
a = 8'd215; b = 8'd123;  #10 
a = 8'd215; b = 8'd124;  #10 
a = 8'd215; b = 8'd125;  #10 
a = 8'd215; b = 8'd126;  #10 
a = 8'd215; b = 8'd127;  #10 
a = 8'd215; b = 8'd128;  #10 
a = 8'd215; b = 8'd129;  #10 
a = 8'd215; b = 8'd130;  #10 
a = 8'd215; b = 8'd131;  #10 
a = 8'd215; b = 8'd132;  #10 
a = 8'd215; b = 8'd133;  #10 
a = 8'd215; b = 8'd134;  #10 
a = 8'd215; b = 8'd135;  #10 
a = 8'd215; b = 8'd136;  #10 
a = 8'd215; b = 8'd137;  #10 
a = 8'd215; b = 8'd138;  #10 
a = 8'd215; b = 8'd139;  #10 
a = 8'd215; b = 8'd140;  #10 
a = 8'd215; b = 8'd141;  #10 
a = 8'd215; b = 8'd142;  #10 
a = 8'd215; b = 8'd143;  #10 
a = 8'd215; b = 8'd144;  #10 
a = 8'd215; b = 8'd145;  #10 
a = 8'd215; b = 8'd146;  #10 
a = 8'd215; b = 8'd147;  #10 
a = 8'd215; b = 8'd148;  #10 
a = 8'd215; b = 8'd149;  #10 
a = 8'd215; b = 8'd150;  #10 
a = 8'd215; b = 8'd151;  #10 
a = 8'd215; b = 8'd152;  #10 
a = 8'd215; b = 8'd153;  #10 
a = 8'd215; b = 8'd154;  #10 
a = 8'd215; b = 8'd155;  #10 
a = 8'd215; b = 8'd156;  #10 
a = 8'd215; b = 8'd157;  #10 
a = 8'd215; b = 8'd158;  #10 
a = 8'd215; b = 8'd159;  #10 
a = 8'd215; b = 8'd160;  #10 
a = 8'd215; b = 8'd161;  #10 
a = 8'd215; b = 8'd162;  #10 
a = 8'd215; b = 8'd163;  #10 
a = 8'd215; b = 8'd164;  #10 
a = 8'd215; b = 8'd165;  #10 
a = 8'd215; b = 8'd166;  #10 
a = 8'd215; b = 8'd167;  #10 
a = 8'd215; b = 8'd168;  #10 
a = 8'd215; b = 8'd169;  #10 
a = 8'd215; b = 8'd170;  #10 
a = 8'd215; b = 8'd171;  #10 
a = 8'd215; b = 8'd172;  #10 
a = 8'd215; b = 8'd173;  #10 
a = 8'd215; b = 8'd174;  #10 
a = 8'd215; b = 8'd175;  #10 
a = 8'd215; b = 8'd176;  #10 
a = 8'd215; b = 8'd177;  #10 
a = 8'd215; b = 8'd178;  #10 
a = 8'd215; b = 8'd179;  #10 
a = 8'd215; b = 8'd180;  #10 
a = 8'd215; b = 8'd181;  #10 
a = 8'd215; b = 8'd182;  #10 
a = 8'd215; b = 8'd183;  #10 
a = 8'd215; b = 8'd184;  #10 
a = 8'd215; b = 8'd185;  #10 
a = 8'd215; b = 8'd186;  #10 
a = 8'd215; b = 8'd187;  #10 
a = 8'd215; b = 8'd188;  #10 
a = 8'd215; b = 8'd189;  #10 
a = 8'd215; b = 8'd190;  #10 
a = 8'd215; b = 8'd191;  #10 
a = 8'd215; b = 8'd192;  #10 
a = 8'd215; b = 8'd193;  #10 
a = 8'd215; b = 8'd194;  #10 
a = 8'd215; b = 8'd195;  #10 
a = 8'd215; b = 8'd196;  #10 
a = 8'd215; b = 8'd197;  #10 
a = 8'd215; b = 8'd198;  #10 
a = 8'd215; b = 8'd199;  #10 
a = 8'd215; b = 8'd200;  #10 
a = 8'd215; b = 8'd201;  #10 
a = 8'd215; b = 8'd202;  #10 
a = 8'd215; b = 8'd203;  #10 
a = 8'd215; b = 8'd204;  #10 
a = 8'd215; b = 8'd205;  #10 
a = 8'd215; b = 8'd206;  #10 
a = 8'd215; b = 8'd207;  #10 
a = 8'd215; b = 8'd208;  #10 
a = 8'd215; b = 8'd209;  #10 
a = 8'd215; b = 8'd210;  #10 
a = 8'd215; b = 8'd211;  #10 
a = 8'd215; b = 8'd212;  #10 
a = 8'd215; b = 8'd213;  #10 
a = 8'd215; b = 8'd214;  #10 
a = 8'd215; b = 8'd215;  #10 
a = 8'd215; b = 8'd216;  #10 
a = 8'd215; b = 8'd217;  #10 
a = 8'd215; b = 8'd218;  #10 
a = 8'd215; b = 8'd219;  #10 
a = 8'd215; b = 8'd220;  #10 
a = 8'd215; b = 8'd221;  #10 
a = 8'd215; b = 8'd222;  #10 
a = 8'd215; b = 8'd223;  #10 
a = 8'd215; b = 8'd224;  #10 
a = 8'd215; b = 8'd225;  #10 
a = 8'd215; b = 8'd226;  #10 
a = 8'd215; b = 8'd227;  #10 
a = 8'd215; b = 8'd228;  #10 
a = 8'd215; b = 8'd229;  #10 
a = 8'd215; b = 8'd230;  #10 
a = 8'd215; b = 8'd231;  #10 
a = 8'd215; b = 8'd232;  #10 
a = 8'd215; b = 8'd233;  #10 
a = 8'd215; b = 8'd234;  #10 
a = 8'd215; b = 8'd235;  #10 
a = 8'd215; b = 8'd236;  #10 
a = 8'd215; b = 8'd237;  #10 
a = 8'd215; b = 8'd238;  #10 
a = 8'd215; b = 8'd239;  #10 
a = 8'd215; b = 8'd240;  #10 
a = 8'd215; b = 8'd241;  #10 
a = 8'd215; b = 8'd242;  #10 
a = 8'd215; b = 8'd243;  #10 
a = 8'd215; b = 8'd244;  #10 
a = 8'd215; b = 8'd245;  #10 
a = 8'd215; b = 8'd246;  #10 
a = 8'd215; b = 8'd247;  #10 
a = 8'd215; b = 8'd248;  #10 
a = 8'd215; b = 8'd249;  #10 
a = 8'd215; b = 8'd250;  #10 
a = 8'd215; b = 8'd251;  #10 
a = 8'd215; b = 8'd252;  #10 
a = 8'd215; b = 8'd253;  #10 
a = 8'd215; b = 8'd254;  #10 
a = 8'd215; b = 8'd255;  #10 
a = 8'd216; b = 8'd0;  #10 
a = 8'd216; b = 8'd1;  #10 
a = 8'd216; b = 8'd2;  #10 
a = 8'd216; b = 8'd3;  #10 
a = 8'd216; b = 8'd4;  #10 
a = 8'd216; b = 8'd5;  #10 
a = 8'd216; b = 8'd6;  #10 
a = 8'd216; b = 8'd7;  #10 
a = 8'd216; b = 8'd8;  #10 
a = 8'd216; b = 8'd9;  #10 
a = 8'd216; b = 8'd10;  #10 
a = 8'd216; b = 8'd11;  #10 
a = 8'd216; b = 8'd12;  #10 
a = 8'd216; b = 8'd13;  #10 
a = 8'd216; b = 8'd14;  #10 
a = 8'd216; b = 8'd15;  #10 
a = 8'd216; b = 8'd16;  #10 
a = 8'd216; b = 8'd17;  #10 
a = 8'd216; b = 8'd18;  #10 
a = 8'd216; b = 8'd19;  #10 
a = 8'd216; b = 8'd20;  #10 
a = 8'd216; b = 8'd21;  #10 
a = 8'd216; b = 8'd22;  #10 
a = 8'd216; b = 8'd23;  #10 
a = 8'd216; b = 8'd24;  #10 
a = 8'd216; b = 8'd25;  #10 
a = 8'd216; b = 8'd26;  #10 
a = 8'd216; b = 8'd27;  #10 
a = 8'd216; b = 8'd28;  #10 
a = 8'd216; b = 8'd29;  #10 
a = 8'd216; b = 8'd30;  #10 
a = 8'd216; b = 8'd31;  #10 
a = 8'd216; b = 8'd32;  #10 
a = 8'd216; b = 8'd33;  #10 
a = 8'd216; b = 8'd34;  #10 
a = 8'd216; b = 8'd35;  #10 
a = 8'd216; b = 8'd36;  #10 
a = 8'd216; b = 8'd37;  #10 
a = 8'd216; b = 8'd38;  #10 
a = 8'd216; b = 8'd39;  #10 
a = 8'd216; b = 8'd40;  #10 
a = 8'd216; b = 8'd41;  #10 
a = 8'd216; b = 8'd42;  #10 
a = 8'd216; b = 8'd43;  #10 
a = 8'd216; b = 8'd44;  #10 
a = 8'd216; b = 8'd45;  #10 
a = 8'd216; b = 8'd46;  #10 
a = 8'd216; b = 8'd47;  #10 
a = 8'd216; b = 8'd48;  #10 
a = 8'd216; b = 8'd49;  #10 
a = 8'd216; b = 8'd50;  #10 
a = 8'd216; b = 8'd51;  #10 
a = 8'd216; b = 8'd52;  #10 
a = 8'd216; b = 8'd53;  #10 
a = 8'd216; b = 8'd54;  #10 
a = 8'd216; b = 8'd55;  #10 
a = 8'd216; b = 8'd56;  #10 
a = 8'd216; b = 8'd57;  #10 
a = 8'd216; b = 8'd58;  #10 
a = 8'd216; b = 8'd59;  #10 
a = 8'd216; b = 8'd60;  #10 
a = 8'd216; b = 8'd61;  #10 
a = 8'd216; b = 8'd62;  #10 
a = 8'd216; b = 8'd63;  #10 
a = 8'd216; b = 8'd64;  #10 
a = 8'd216; b = 8'd65;  #10 
a = 8'd216; b = 8'd66;  #10 
a = 8'd216; b = 8'd67;  #10 
a = 8'd216; b = 8'd68;  #10 
a = 8'd216; b = 8'd69;  #10 
a = 8'd216; b = 8'd70;  #10 
a = 8'd216; b = 8'd71;  #10 
a = 8'd216; b = 8'd72;  #10 
a = 8'd216; b = 8'd73;  #10 
a = 8'd216; b = 8'd74;  #10 
a = 8'd216; b = 8'd75;  #10 
a = 8'd216; b = 8'd76;  #10 
a = 8'd216; b = 8'd77;  #10 
a = 8'd216; b = 8'd78;  #10 
a = 8'd216; b = 8'd79;  #10 
a = 8'd216; b = 8'd80;  #10 
a = 8'd216; b = 8'd81;  #10 
a = 8'd216; b = 8'd82;  #10 
a = 8'd216; b = 8'd83;  #10 
a = 8'd216; b = 8'd84;  #10 
a = 8'd216; b = 8'd85;  #10 
a = 8'd216; b = 8'd86;  #10 
a = 8'd216; b = 8'd87;  #10 
a = 8'd216; b = 8'd88;  #10 
a = 8'd216; b = 8'd89;  #10 
a = 8'd216; b = 8'd90;  #10 
a = 8'd216; b = 8'd91;  #10 
a = 8'd216; b = 8'd92;  #10 
a = 8'd216; b = 8'd93;  #10 
a = 8'd216; b = 8'd94;  #10 
a = 8'd216; b = 8'd95;  #10 
a = 8'd216; b = 8'd96;  #10 
a = 8'd216; b = 8'd97;  #10 
a = 8'd216; b = 8'd98;  #10 
a = 8'd216; b = 8'd99;  #10 
a = 8'd216; b = 8'd100;  #10 
a = 8'd216; b = 8'd101;  #10 
a = 8'd216; b = 8'd102;  #10 
a = 8'd216; b = 8'd103;  #10 
a = 8'd216; b = 8'd104;  #10 
a = 8'd216; b = 8'd105;  #10 
a = 8'd216; b = 8'd106;  #10 
a = 8'd216; b = 8'd107;  #10 
a = 8'd216; b = 8'd108;  #10 
a = 8'd216; b = 8'd109;  #10 
a = 8'd216; b = 8'd110;  #10 
a = 8'd216; b = 8'd111;  #10 
a = 8'd216; b = 8'd112;  #10 
a = 8'd216; b = 8'd113;  #10 
a = 8'd216; b = 8'd114;  #10 
a = 8'd216; b = 8'd115;  #10 
a = 8'd216; b = 8'd116;  #10 
a = 8'd216; b = 8'd117;  #10 
a = 8'd216; b = 8'd118;  #10 
a = 8'd216; b = 8'd119;  #10 
a = 8'd216; b = 8'd120;  #10 
a = 8'd216; b = 8'd121;  #10 
a = 8'd216; b = 8'd122;  #10 
a = 8'd216; b = 8'd123;  #10 
a = 8'd216; b = 8'd124;  #10 
a = 8'd216; b = 8'd125;  #10 
a = 8'd216; b = 8'd126;  #10 
a = 8'd216; b = 8'd127;  #10 
a = 8'd216; b = 8'd128;  #10 
a = 8'd216; b = 8'd129;  #10 
a = 8'd216; b = 8'd130;  #10 
a = 8'd216; b = 8'd131;  #10 
a = 8'd216; b = 8'd132;  #10 
a = 8'd216; b = 8'd133;  #10 
a = 8'd216; b = 8'd134;  #10 
a = 8'd216; b = 8'd135;  #10 
a = 8'd216; b = 8'd136;  #10 
a = 8'd216; b = 8'd137;  #10 
a = 8'd216; b = 8'd138;  #10 
a = 8'd216; b = 8'd139;  #10 
a = 8'd216; b = 8'd140;  #10 
a = 8'd216; b = 8'd141;  #10 
a = 8'd216; b = 8'd142;  #10 
a = 8'd216; b = 8'd143;  #10 
a = 8'd216; b = 8'd144;  #10 
a = 8'd216; b = 8'd145;  #10 
a = 8'd216; b = 8'd146;  #10 
a = 8'd216; b = 8'd147;  #10 
a = 8'd216; b = 8'd148;  #10 
a = 8'd216; b = 8'd149;  #10 
a = 8'd216; b = 8'd150;  #10 
a = 8'd216; b = 8'd151;  #10 
a = 8'd216; b = 8'd152;  #10 
a = 8'd216; b = 8'd153;  #10 
a = 8'd216; b = 8'd154;  #10 
a = 8'd216; b = 8'd155;  #10 
a = 8'd216; b = 8'd156;  #10 
a = 8'd216; b = 8'd157;  #10 
a = 8'd216; b = 8'd158;  #10 
a = 8'd216; b = 8'd159;  #10 
a = 8'd216; b = 8'd160;  #10 
a = 8'd216; b = 8'd161;  #10 
a = 8'd216; b = 8'd162;  #10 
a = 8'd216; b = 8'd163;  #10 
a = 8'd216; b = 8'd164;  #10 
a = 8'd216; b = 8'd165;  #10 
a = 8'd216; b = 8'd166;  #10 
a = 8'd216; b = 8'd167;  #10 
a = 8'd216; b = 8'd168;  #10 
a = 8'd216; b = 8'd169;  #10 
a = 8'd216; b = 8'd170;  #10 
a = 8'd216; b = 8'd171;  #10 
a = 8'd216; b = 8'd172;  #10 
a = 8'd216; b = 8'd173;  #10 
a = 8'd216; b = 8'd174;  #10 
a = 8'd216; b = 8'd175;  #10 
a = 8'd216; b = 8'd176;  #10 
a = 8'd216; b = 8'd177;  #10 
a = 8'd216; b = 8'd178;  #10 
a = 8'd216; b = 8'd179;  #10 
a = 8'd216; b = 8'd180;  #10 
a = 8'd216; b = 8'd181;  #10 
a = 8'd216; b = 8'd182;  #10 
a = 8'd216; b = 8'd183;  #10 
a = 8'd216; b = 8'd184;  #10 
a = 8'd216; b = 8'd185;  #10 
a = 8'd216; b = 8'd186;  #10 
a = 8'd216; b = 8'd187;  #10 
a = 8'd216; b = 8'd188;  #10 
a = 8'd216; b = 8'd189;  #10 
a = 8'd216; b = 8'd190;  #10 
a = 8'd216; b = 8'd191;  #10 
a = 8'd216; b = 8'd192;  #10 
a = 8'd216; b = 8'd193;  #10 
a = 8'd216; b = 8'd194;  #10 
a = 8'd216; b = 8'd195;  #10 
a = 8'd216; b = 8'd196;  #10 
a = 8'd216; b = 8'd197;  #10 
a = 8'd216; b = 8'd198;  #10 
a = 8'd216; b = 8'd199;  #10 
a = 8'd216; b = 8'd200;  #10 
a = 8'd216; b = 8'd201;  #10 
a = 8'd216; b = 8'd202;  #10 
a = 8'd216; b = 8'd203;  #10 
a = 8'd216; b = 8'd204;  #10 
a = 8'd216; b = 8'd205;  #10 
a = 8'd216; b = 8'd206;  #10 
a = 8'd216; b = 8'd207;  #10 
a = 8'd216; b = 8'd208;  #10 
a = 8'd216; b = 8'd209;  #10 
a = 8'd216; b = 8'd210;  #10 
a = 8'd216; b = 8'd211;  #10 
a = 8'd216; b = 8'd212;  #10 
a = 8'd216; b = 8'd213;  #10 
a = 8'd216; b = 8'd214;  #10 
a = 8'd216; b = 8'd215;  #10 
a = 8'd216; b = 8'd216;  #10 
a = 8'd216; b = 8'd217;  #10 
a = 8'd216; b = 8'd218;  #10 
a = 8'd216; b = 8'd219;  #10 
a = 8'd216; b = 8'd220;  #10 
a = 8'd216; b = 8'd221;  #10 
a = 8'd216; b = 8'd222;  #10 
a = 8'd216; b = 8'd223;  #10 
a = 8'd216; b = 8'd224;  #10 
a = 8'd216; b = 8'd225;  #10 
a = 8'd216; b = 8'd226;  #10 
a = 8'd216; b = 8'd227;  #10 
a = 8'd216; b = 8'd228;  #10 
a = 8'd216; b = 8'd229;  #10 
a = 8'd216; b = 8'd230;  #10 
a = 8'd216; b = 8'd231;  #10 
a = 8'd216; b = 8'd232;  #10 
a = 8'd216; b = 8'd233;  #10 
a = 8'd216; b = 8'd234;  #10 
a = 8'd216; b = 8'd235;  #10 
a = 8'd216; b = 8'd236;  #10 
a = 8'd216; b = 8'd237;  #10 
a = 8'd216; b = 8'd238;  #10 
a = 8'd216; b = 8'd239;  #10 
a = 8'd216; b = 8'd240;  #10 
a = 8'd216; b = 8'd241;  #10 
a = 8'd216; b = 8'd242;  #10 
a = 8'd216; b = 8'd243;  #10 
a = 8'd216; b = 8'd244;  #10 
a = 8'd216; b = 8'd245;  #10 
a = 8'd216; b = 8'd246;  #10 
a = 8'd216; b = 8'd247;  #10 
a = 8'd216; b = 8'd248;  #10 
a = 8'd216; b = 8'd249;  #10 
a = 8'd216; b = 8'd250;  #10 
a = 8'd216; b = 8'd251;  #10 
a = 8'd216; b = 8'd252;  #10 
a = 8'd216; b = 8'd253;  #10 
a = 8'd216; b = 8'd254;  #10 
a = 8'd216; b = 8'd255;  #10 
a = 8'd217; b = 8'd0;  #10 
a = 8'd217; b = 8'd1;  #10 
a = 8'd217; b = 8'd2;  #10 
a = 8'd217; b = 8'd3;  #10 
a = 8'd217; b = 8'd4;  #10 
a = 8'd217; b = 8'd5;  #10 
a = 8'd217; b = 8'd6;  #10 
a = 8'd217; b = 8'd7;  #10 
a = 8'd217; b = 8'd8;  #10 
a = 8'd217; b = 8'd9;  #10 
a = 8'd217; b = 8'd10;  #10 
a = 8'd217; b = 8'd11;  #10 
a = 8'd217; b = 8'd12;  #10 
a = 8'd217; b = 8'd13;  #10 
a = 8'd217; b = 8'd14;  #10 
a = 8'd217; b = 8'd15;  #10 
a = 8'd217; b = 8'd16;  #10 
a = 8'd217; b = 8'd17;  #10 
a = 8'd217; b = 8'd18;  #10 
a = 8'd217; b = 8'd19;  #10 
a = 8'd217; b = 8'd20;  #10 
a = 8'd217; b = 8'd21;  #10 
a = 8'd217; b = 8'd22;  #10 
a = 8'd217; b = 8'd23;  #10 
a = 8'd217; b = 8'd24;  #10 
a = 8'd217; b = 8'd25;  #10 
a = 8'd217; b = 8'd26;  #10 
a = 8'd217; b = 8'd27;  #10 
a = 8'd217; b = 8'd28;  #10 
a = 8'd217; b = 8'd29;  #10 
a = 8'd217; b = 8'd30;  #10 
a = 8'd217; b = 8'd31;  #10 
a = 8'd217; b = 8'd32;  #10 
a = 8'd217; b = 8'd33;  #10 
a = 8'd217; b = 8'd34;  #10 
a = 8'd217; b = 8'd35;  #10 
a = 8'd217; b = 8'd36;  #10 
a = 8'd217; b = 8'd37;  #10 
a = 8'd217; b = 8'd38;  #10 
a = 8'd217; b = 8'd39;  #10 
a = 8'd217; b = 8'd40;  #10 
a = 8'd217; b = 8'd41;  #10 
a = 8'd217; b = 8'd42;  #10 
a = 8'd217; b = 8'd43;  #10 
a = 8'd217; b = 8'd44;  #10 
a = 8'd217; b = 8'd45;  #10 
a = 8'd217; b = 8'd46;  #10 
a = 8'd217; b = 8'd47;  #10 
a = 8'd217; b = 8'd48;  #10 
a = 8'd217; b = 8'd49;  #10 
a = 8'd217; b = 8'd50;  #10 
a = 8'd217; b = 8'd51;  #10 
a = 8'd217; b = 8'd52;  #10 
a = 8'd217; b = 8'd53;  #10 
a = 8'd217; b = 8'd54;  #10 
a = 8'd217; b = 8'd55;  #10 
a = 8'd217; b = 8'd56;  #10 
a = 8'd217; b = 8'd57;  #10 
a = 8'd217; b = 8'd58;  #10 
a = 8'd217; b = 8'd59;  #10 
a = 8'd217; b = 8'd60;  #10 
a = 8'd217; b = 8'd61;  #10 
a = 8'd217; b = 8'd62;  #10 
a = 8'd217; b = 8'd63;  #10 
a = 8'd217; b = 8'd64;  #10 
a = 8'd217; b = 8'd65;  #10 
a = 8'd217; b = 8'd66;  #10 
a = 8'd217; b = 8'd67;  #10 
a = 8'd217; b = 8'd68;  #10 
a = 8'd217; b = 8'd69;  #10 
a = 8'd217; b = 8'd70;  #10 
a = 8'd217; b = 8'd71;  #10 
a = 8'd217; b = 8'd72;  #10 
a = 8'd217; b = 8'd73;  #10 
a = 8'd217; b = 8'd74;  #10 
a = 8'd217; b = 8'd75;  #10 
a = 8'd217; b = 8'd76;  #10 
a = 8'd217; b = 8'd77;  #10 
a = 8'd217; b = 8'd78;  #10 
a = 8'd217; b = 8'd79;  #10 
a = 8'd217; b = 8'd80;  #10 
a = 8'd217; b = 8'd81;  #10 
a = 8'd217; b = 8'd82;  #10 
a = 8'd217; b = 8'd83;  #10 
a = 8'd217; b = 8'd84;  #10 
a = 8'd217; b = 8'd85;  #10 
a = 8'd217; b = 8'd86;  #10 
a = 8'd217; b = 8'd87;  #10 
a = 8'd217; b = 8'd88;  #10 
a = 8'd217; b = 8'd89;  #10 
a = 8'd217; b = 8'd90;  #10 
a = 8'd217; b = 8'd91;  #10 
a = 8'd217; b = 8'd92;  #10 
a = 8'd217; b = 8'd93;  #10 
a = 8'd217; b = 8'd94;  #10 
a = 8'd217; b = 8'd95;  #10 
a = 8'd217; b = 8'd96;  #10 
a = 8'd217; b = 8'd97;  #10 
a = 8'd217; b = 8'd98;  #10 
a = 8'd217; b = 8'd99;  #10 
a = 8'd217; b = 8'd100;  #10 
a = 8'd217; b = 8'd101;  #10 
a = 8'd217; b = 8'd102;  #10 
a = 8'd217; b = 8'd103;  #10 
a = 8'd217; b = 8'd104;  #10 
a = 8'd217; b = 8'd105;  #10 
a = 8'd217; b = 8'd106;  #10 
a = 8'd217; b = 8'd107;  #10 
a = 8'd217; b = 8'd108;  #10 
a = 8'd217; b = 8'd109;  #10 
a = 8'd217; b = 8'd110;  #10 
a = 8'd217; b = 8'd111;  #10 
a = 8'd217; b = 8'd112;  #10 
a = 8'd217; b = 8'd113;  #10 
a = 8'd217; b = 8'd114;  #10 
a = 8'd217; b = 8'd115;  #10 
a = 8'd217; b = 8'd116;  #10 
a = 8'd217; b = 8'd117;  #10 
a = 8'd217; b = 8'd118;  #10 
a = 8'd217; b = 8'd119;  #10 
a = 8'd217; b = 8'd120;  #10 
a = 8'd217; b = 8'd121;  #10 
a = 8'd217; b = 8'd122;  #10 
a = 8'd217; b = 8'd123;  #10 
a = 8'd217; b = 8'd124;  #10 
a = 8'd217; b = 8'd125;  #10 
a = 8'd217; b = 8'd126;  #10 
a = 8'd217; b = 8'd127;  #10 
a = 8'd217; b = 8'd128;  #10 
a = 8'd217; b = 8'd129;  #10 
a = 8'd217; b = 8'd130;  #10 
a = 8'd217; b = 8'd131;  #10 
a = 8'd217; b = 8'd132;  #10 
a = 8'd217; b = 8'd133;  #10 
a = 8'd217; b = 8'd134;  #10 
a = 8'd217; b = 8'd135;  #10 
a = 8'd217; b = 8'd136;  #10 
a = 8'd217; b = 8'd137;  #10 
a = 8'd217; b = 8'd138;  #10 
a = 8'd217; b = 8'd139;  #10 
a = 8'd217; b = 8'd140;  #10 
a = 8'd217; b = 8'd141;  #10 
a = 8'd217; b = 8'd142;  #10 
a = 8'd217; b = 8'd143;  #10 
a = 8'd217; b = 8'd144;  #10 
a = 8'd217; b = 8'd145;  #10 
a = 8'd217; b = 8'd146;  #10 
a = 8'd217; b = 8'd147;  #10 
a = 8'd217; b = 8'd148;  #10 
a = 8'd217; b = 8'd149;  #10 
a = 8'd217; b = 8'd150;  #10 
a = 8'd217; b = 8'd151;  #10 
a = 8'd217; b = 8'd152;  #10 
a = 8'd217; b = 8'd153;  #10 
a = 8'd217; b = 8'd154;  #10 
a = 8'd217; b = 8'd155;  #10 
a = 8'd217; b = 8'd156;  #10 
a = 8'd217; b = 8'd157;  #10 
a = 8'd217; b = 8'd158;  #10 
a = 8'd217; b = 8'd159;  #10 
a = 8'd217; b = 8'd160;  #10 
a = 8'd217; b = 8'd161;  #10 
a = 8'd217; b = 8'd162;  #10 
a = 8'd217; b = 8'd163;  #10 
a = 8'd217; b = 8'd164;  #10 
a = 8'd217; b = 8'd165;  #10 
a = 8'd217; b = 8'd166;  #10 
a = 8'd217; b = 8'd167;  #10 
a = 8'd217; b = 8'd168;  #10 
a = 8'd217; b = 8'd169;  #10 
a = 8'd217; b = 8'd170;  #10 
a = 8'd217; b = 8'd171;  #10 
a = 8'd217; b = 8'd172;  #10 
a = 8'd217; b = 8'd173;  #10 
a = 8'd217; b = 8'd174;  #10 
a = 8'd217; b = 8'd175;  #10 
a = 8'd217; b = 8'd176;  #10 
a = 8'd217; b = 8'd177;  #10 
a = 8'd217; b = 8'd178;  #10 
a = 8'd217; b = 8'd179;  #10 
a = 8'd217; b = 8'd180;  #10 
a = 8'd217; b = 8'd181;  #10 
a = 8'd217; b = 8'd182;  #10 
a = 8'd217; b = 8'd183;  #10 
a = 8'd217; b = 8'd184;  #10 
a = 8'd217; b = 8'd185;  #10 
a = 8'd217; b = 8'd186;  #10 
a = 8'd217; b = 8'd187;  #10 
a = 8'd217; b = 8'd188;  #10 
a = 8'd217; b = 8'd189;  #10 
a = 8'd217; b = 8'd190;  #10 
a = 8'd217; b = 8'd191;  #10 
a = 8'd217; b = 8'd192;  #10 
a = 8'd217; b = 8'd193;  #10 
a = 8'd217; b = 8'd194;  #10 
a = 8'd217; b = 8'd195;  #10 
a = 8'd217; b = 8'd196;  #10 
a = 8'd217; b = 8'd197;  #10 
a = 8'd217; b = 8'd198;  #10 
a = 8'd217; b = 8'd199;  #10 
a = 8'd217; b = 8'd200;  #10 
a = 8'd217; b = 8'd201;  #10 
a = 8'd217; b = 8'd202;  #10 
a = 8'd217; b = 8'd203;  #10 
a = 8'd217; b = 8'd204;  #10 
a = 8'd217; b = 8'd205;  #10 
a = 8'd217; b = 8'd206;  #10 
a = 8'd217; b = 8'd207;  #10 
a = 8'd217; b = 8'd208;  #10 
a = 8'd217; b = 8'd209;  #10 
a = 8'd217; b = 8'd210;  #10 
a = 8'd217; b = 8'd211;  #10 
a = 8'd217; b = 8'd212;  #10 
a = 8'd217; b = 8'd213;  #10 
a = 8'd217; b = 8'd214;  #10 
a = 8'd217; b = 8'd215;  #10 
a = 8'd217; b = 8'd216;  #10 
a = 8'd217; b = 8'd217;  #10 
a = 8'd217; b = 8'd218;  #10 
a = 8'd217; b = 8'd219;  #10 
a = 8'd217; b = 8'd220;  #10 
a = 8'd217; b = 8'd221;  #10 
a = 8'd217; b = 8'd222;  #10 
a = 8'd217; b = 8'd223;  #10 
a = 8'd217; b = 8'd224;  #10 
a = 8'd217; b = 8'd225;  #10 
a = 8'd217; b = 8'd226;  #10 
a = 8'd217; b = 8'd227;  #10 
a = 8'd217; b = 8'd228;  #10 
a = 8'd217; b = 8'd229;  #10 
a = 8'd217; b = 8'd230;  #10 
a = 8'd217; b = 8'd231;  #10 
a = 8'd217; b = 8'd232;  #10 
a = 8'd217; b = 8'd233;  #10 
a = 8'd217; b = 8'd234;  #10 
a = 8'd217; b = 8'd235;  #10 
a = 8'd217; b = 8'd236;  #10 
a = 8'd217; b = 8'd237;  #10 
a = 8'd217; b = 8'd238;  #10 
a = 8'd217; b = 8'd239;  #10 
a = 8'd217; b = 8'd240;  #10 
a = 8'd217; b = 8'd241;  #10 
a = 8'd217; b = 8'd242;  #10 
a = 8'd217; b = 8'd243;  #10 
a = 8'd217; b = 8'd244;  #10 
a = 8'd217; b = 8'd245;  #10 
a = 8'd217; b = 8'd246;  #10 
a = 8'd217; b = 8'd247;  #10 
a = 8'd217; b = 8'd248;  #10 
a = 8'd217; b = 8'd249;  #10 
a = 8'd217; b = 8'd250;  #10 
a = 8'd217; b = 8'd251;  #10 
a = 8'd217; b = 8'd252;  #10 
a = 8'd217; b = 8'd253;  #10 
a = 8'd217; b = 8'd254;  #10 
a = 8'd217; b = 8'd255;  #10 
a = 8'd218; b = 8'd0;  #10 
a = 8'd218; b = 8'd1;  #10 
a = 8'd218; b = 8'd2;  #10 
a = 8'd218; b = 8'd3;  #10 
a = 8'd218; b = 8'd4;  #10 
a = 8'd218; b = 8'd5;  #10 
a = 8'd218; b = 8'd6;  #10 
a = 8'd218; b = 8'd7;  #10 
a = 8'd218; b = 8'd8;  #10 
a = 8'd218; b = 8'd9;  #10 
a = 8'd218; b = 8'd10;  #10 
a = 8'd218; b = 8'd11;  #10 
a = 8'd218; b = 8'd12;  #10 
a = 8'd218; b = 8'd13;  #10 
a = 8'd218; b = 8'd14;  #10 
a = 8'd218; b = 8'd15;  #10 
a = 8'd218; b = 8'd16;  #10 
a = 8'd218; b = 8'd17;  #10 
a = 8'd218; b = 8'd18;  #10 
a = 8'd218; b = 8'd19;  #10 
a = 8'd218; b = 8'd20;  #10 
a = 8'd218; b = 8'd21;  #10 
a = 8'd218; b = 8'd22;  #10 
a = 8'd218; b = 8'd23;  #10 
a = 8'd218; b = 8'd24;  #10 
a = 8'd218; b = 8'd25;  #10 
a = 8'd218; b = 8'd26;  #10 
a = 8'd218; b = 8'd27;  #10 
a = 8'd218; b = 8'd28;  #10 
a = 8'd218; b = 8'd29;  #10 
a = 8'd218; b = 8'd30;  #10 
a = 8'd218; b = 8'd31;  #10 
a = 8'd218; b = 8'd32;  #10 
a = 8'd218; b = 8'd33;  #10 
a = 8'd218; b = 8'd34;  #10 
a = 8'd218; b = 8'd35;  #10 
a = 8'd218; b = 8'd36;  #10 
a = 8'd218; b = 8'd37;  #10 
a = 8'd218; b = 8'd38;  #10 
a = 8'd218; b = 8'd39;  #10 
a = 8'd218; b = 8'd40;  #10 
a = 8'd218; b = 8'd41;  #10 
a = 8'd218; b = 8'd42;  #10 
a = 8'd218; b = 8'd43;  #10 
a = 8'd218; b = 8'd44;  #10 
a = 8'd218; b = 8'd45;  #10 
a = 8'd218; b = 8'd46;  #10 
a = 8'd218; b = 8'd47;  #10 
a = 8'd218; b = 8'd48;  #10 
a = 8'd218; b = 8'd49;  #10 
a = 8'd218; b = 8'd50;  #10 
a = 8'd218; b = 8'd51;  #10 
a = 8'd218; b = 8'd52;  #10 
a = 8'd218; b = 8'd53;  #10 
a = 8'd218; b = 8'd54;  #10 
a = 8'd218; b = 8'd55;  #10 
a = 8'd218; b = 8'd56;  #10 
a = 8'd218; b = 8'd57;  #10 
a = 8'd218; b = 8'd58;  #10 
a = 8'd218; b = 8'd59;  #10 
a = 8'd218; b = 8'd60;  #10 
a = 8'd218; b = 8'd61;  #10 
a = 8'd218; b = 8'd62;  #10 
a = 8'd218; b = 8'd63;  #10 
a = 8'd218; b = 8'd64;  #10 
a = 8'd218; b = 8'd65;  #10 
a = 8'd218; b = 8'd66;  #10 
a = 8'd218; b = 8'd67;  #10 
a = 8'd218; b = 8'd68;  #10 
a = 8'd218; b = 8'd69;  #10 
a = 8'd218; b = 8'd70;  #10 
a = 8'd218; b = 8'd71;  #10 
a = 8'd218; b = 8'd72;  #10 
a = 8'd218; b = 8'd73;  #10 
a = 8'd218; b = 8'd74;  #10 
a = 8'd218; b = 8'd75;  #10 
a = 8'd218; b = 8'd76;  #10 
a = 8'd218; b = 8'd77;  #10 
a = 8'd218; b = 8'd78;  #10 
a = 8'd218; b = 8'd79;  #10 
a = 8'd218; b = 8'd80;  #10 
a = 8'd218; b = 8'd81;  #10 
a = 8'd218; b = 8'd82;  #10 
a = 8'd218; b = 8'd83;  #10 
a = 8'd218; b = 8'd84;  #10 
a = 8'd218; b = 8'd85;  #10 
a = 8'd218; b = 8'd86;  #10 
a = 8'd218; b = 8'd87;  #10 
a = 8'd218; b = 8'd88;  #10 
a = 8'd218; b = 8'd89;  #10 
a = 8'd218; b = 8'd90;  #10 
a = 8'd218; b = 8'd91;  #10 
a = 8'd218; b = 8'd92;  #10 
a = 8'd218; b = 8'd93;  #10 
a = 8'd218; b = 8'd94;  #10 
a = 8'd218; b = 8'd95;  #10 
a = 8'd218; b = 8'd96;  #10 
a = 8'd218; b = 8'd97;  #10 
a = 8'd218; b = 8'd98;  #10 
a = 8'd218; b = 8'd99;  #10 
a = 8'd218; b = 8'd100;  #10 
a = 8'd218; b = 8'd101;  #10 
a = 8'd218; b = 8'd102;  #10 
a = 8'd218; b = 8'd103;  #10 
a = 8'd218; b = 8'd104;  #10 
a = 8'd218; b = 8'd105;  #10 
a = 8'd218; b = 8'd106;  #10 
a = 8'd218; b = 8'd107;  #10 
a = 8'd218; b = 8'd108;  #10 
a = 8'd218; b = 8'd109;  #10 
a = 8'd218; b = 8'd110;  #10 
a = 8'd218; b = 8'd111;  #10 
a = 8'd218; b = 8'd112;  #10 
a = 8'd218; b = 8'd113;  #10 
a = 8'd218; b = 8'd114;  #10 
a = 8'd218; b = 8'd115;  #10 
a = 8'd218; b = 8'd116;  #10 
a = 8'd218; b = 8'd117;  #10 
a = 8'd218; b = 8'd118;  #10 
a = 8'd218; b = 8'd119;  #10 
a = 8'd218; b = 8'd120;  #10 
a = 8'd218; b = 8'd121;  #10 
a = 8'd218; b = 8'd122;  #10 
a = 8'd218; b = 8'd123;  #10 
a = 8'd218; b = 8'd124;  #10 
a = 8'd218; b = 8'd125;  #10 
a = 8'd218; b = 8'd126;  #10 
a = 8'd218; b = 8'd127;  #10 
a = 8'd218; b = 8'd128;  #10 
a = 8'd218; b = 8'd129;  #10 
a = 8'd218; b = 8'd130;  #10 
a = 8'd218; b = 8'd131;  #10 
a = 8'd218; b = 8'd132;  #10 
a = 8'd218; b = 8'd133;  #10 
a = 8'd218; b = 8'd134;  #10 
a = 8'd218; b = 8'd135;  #10 
a = 8'd218; b = 8'd136;  #10 
a = 8'd218; b = 8'd137;  #10 
a = 8'd218; b = 8'd138;  #10 
a = 8'd218; b = 8'd139;  #10 
a = 8'd218; b = 8'd140;  #10 
a = 8'd218; b = 8'd141;  #10 
a = 8'd218; b = 8'd142;  #10 
a = 8'd218; b = 8'd143;  #10 
a = 8'd218; b = 8'd144;  #10 
a = 8'd218; b = 8'd145;  #10 
a = 8'd218; b = 8'd146;  #10 
a = 8'd218; b = 8'd147;  #10 
a = 8'd218; b = 8'd148;  #10 
a = 8'd218; b = 8'd149;  #10 
a = 8'd218; b = 8'd150;  #10 
a = 8'd218; b = 8'd151;  #10 
a = 8'd218; b = 8'd152;  #10 
a = 8'd218; b = 8'd153;  #10 
a = 8'd218; b = 8'd154;  #10 
a = 8'd218; b = 8'd155;  #10 
a = 8'd218; b = 8'd156;  #10 
a = 8'd218; b = 8'd157;  #10 
a = 8'd218; b = 8'd158;  #10 
a = 8'd218; b = 8'd159;  #10 
a = 8'd218; b = 8'd160;  #10 
a = 8'd218; b = 8'd161;  #10 
a = 8'd218; b = 8'd162;  #10 
a = 8'd218; b = 8'd163;  #10 
a = 8'd218; b = 8'd164;  #10 
a = 8'd218; b = 8'd165;  #10 
a = 8'd218; b = 8'd166;  #10 
a = 8'd218; b = 8'd167;  #10 
a = 8'd218; b = 8'd168;  #10 
a = 8'd218; b = 8'd169;  #10 
a = 8'd218; b = 8'd170;  #10 
a = 8'd218; b = 8'd171;  #10 
a = 8'd218; b = 8'd172;  #10 
a = 8'd218; b = 8'd173;  #10 
a = 8'd218; b = 8'd174;  #10 
a = 8'd218; b = 8'd175;  #10 
a = 8'd218; b = 8'd176;  #10 
a = 8'd218; b = 8'd177;  #10 
a = 8'd218; b = 8'd178;  #10 
a = 8'd218; b = 8'd179;  #10 
a = 8'd218; b = 8'd180;  #10 
a = 8'd218; b = 8'd181;  #10 
a = 8'd218; b = 8'd182;  #10 
a = 8'd218; b = 8'd183;  #10 
a = 8'd218; b = 8'd184;  #10 
a = 8'd218; b = 8'd185;  #10 
a = 8'd218; b = 8'd186;  #10 
a = 8'd218; b = 8'd187;  #10 
a = 8'd218; b = 8'd188;  #10 
a = 8'd218; b = 8'd189;  #10 
a = 8'd218; b = 8'd190;  #10 
a = 8'd218; b = 8'd191;  #10 
a = 8'd218; b = 8'd192;  #10 
a = 8'd218; b = 8'd193;  #10 
a = 8'd218; b = 8'd194;  #10 
a = 8'd218; b = 8'd195;  #10 
a = 8'd218; b = 8'd196;  #10 
a = 8'd218; b = 8'd197;  #10 
a = 8'd218; b = 8'd198;  #10 
a = 8'd218; b = 8'd199;  #10 
a = 8'd218; b = 8'd200;  #10 
a = 8'd218; b = 8'd201;  #10 
a = 8'd218; b = 8'd202;  #10 
a = 8'd218; b = 8'd203;  #10 
a = 8'd218; b = 8'd204;  #10 
a = 8'd218; b = 8'd205;  #10 
a = 8'd218; b = 8'd206;  #10 
a = 8'd218; b = 8'd207;  #10 
a = 8'd218; b = 8'd208;  #10 
a = 8'd218; b = 8'd209;  #10 
a = 8'd218; b = 8'd210;  #10 
a = 8'd218; b = 8'd211;  #10 
a = 8'd218; b = 8'd212;  #10 
a = 8'd218; b = 8'd213;  #10 
a = 8'd218; b = 8'd214;  #10 
a = 8'd218; b = 8'd215;  #10 
a = 8'd218; b = 8'd216;  #10 
a = 8'd218; b = 8'd217;  #10 
a = 8'd218; b = 8'd218;  #10 
a = 8'd218; b = 8'd219;  #10 
a = 8'd218; b = 8'd220;  #10 
a = 8'd218; b = 8'd221;  #10 
a = 8'd218; b = 8'd222;  #10 
a = 8'd218; b = 8'd223;  #10 
a = 8'd218; b = 8'd224;  #10 
a = 8'd218; b = 8'd225;  #10 
a = 8'd218; b = 8'd226;  #10 
a = 8'd218; b = 8'd227;  #10 
a = 8'd218; b = 8'd228;  #10 
a = 8'd218; b = 8'd229;  #10 
a = 8'd218; b = 8'd230;  #10 
a = 8'd218; b = 8'd231;  #10 
a = 8'd218; b = 8'd232;  #10 
a = 8'd218; b = 8'd233;  #10 
a = 8'd218; b = 8'd234;  #10 
a = 8'd218; b = 8'd235;  #10 
a = 8'd218; b = 8'd236;  #10 
a = 8'd218; b = 8'd237;  #10 
a = 8'd218; b = 8'd238;  #10 
a = 8'd218; b = 8'd239;  #10 
a = 8'd218; b = 8'd240;  #10 
a = 8'd218; b = 8'd241;  #10 
a = 8'd218; b = 8'd242;  #10 
a = 8'd218; b = 8'd243;  #10 
a = 8'd218; b = 8'd244;  #10 
a = 8'd218; b = 8'd245;  #10 
a = 8'd218; b = 8'd246;  #10 
a = 8'd218; b = 8'd247;  #10 
a = 8'd218; b = 8'd248;  #10 
a = 8'd218; b = 8'd249;  #10 
a = 8'd218; b = 8'd250;  #10 
a = 8'd218; b = 8'd251;  #10 
a = 8'd218; b = 8'd252;  #10 
a = 8'd218; b = 8'd253;  #10 
a = 8'd218; b = 8'd254;  #10 
a = 8'd218; b = 8'd255;  #10 
a = 8'd219; b = 8'd0;  #10 
a = 8'd219; b = 8'd1;  #10 
a = 8'd219; b = 8'd2;  #10 
a = 8'd219; b = 8'd3;  #10 
a = 8'd219; b = 8'd4;  #10 
a = 8'd219; b = 8'd5;  #10 
a = 8'd219; b = 8'd6;  #10 
a = 8'd219; b = 8'd7;  #10 
a = 8'd219; b = 8'd8;  #10 
a = 8'd219; b = 8'd9;  #10 
a = 8'd219; b = 8'd10;  #10 
a = 8'd219; b = 8'd11;  #10 
a = 8'd219; b = 8'd12;  #10 
a = 8'd219; b = 8'd13;  #10 
a = 8'd219; b = 8'd14;  #10 
a = 8'd219; b = 8'd15;  #10 
a = 8'd219; b = 8'd16;  #10 
a = 8'd219; b = 8'd17;  #10 
a = 8'd219; b = 8'd18;  #10 
a = 8'd219; b = 8'd19;  #10 
a = 8'd219; b = 8'd20;  #10 
a = 8'd219; b = 8'd21;  #10 
a = 8'd219; b = 8'd22;  #10 
a = 8'd219; b = 8'd23;  #10 
a = 8'd219; b = 8'd24;  #10 
a = 8'd219; b = 8'd25;  #10 
a = 8'd219; b = 8'd26;  #10 
a = 8'd219; b = 8'd27;  #10 
a = 8'd219; b = 8'd28;  #10 
a = 8'd219; b = 8'd29;  #10 
a = 8'd219; b = 8'd30;  #10 
a = 8'd219; b = 8'd31;  #10 
a = 8'd219; b = 8'd32;  #10 
a = 8'd219; b = 8'd33;  #10 
a = 8'd219; b = 8'd34;  #10 
a = 8'd219; b = 8'd35;  #10 
a = 8'd219; b = 8'd36;  #10 
a = 8'd219; b = 8'd37;  #10 
a = 8'd219; b = 8'd38;  #10 
a = 8'd219; b = 8'd39;  #10 
a = 8'd219; b = 8'd40;  #10 
a = 8'd219; b = 8'd41;  #10 
a = 8'd219; b = 8'd42;  #10 
a = 8'd219; b = 8'd43;  #10 
a = 8'd219; b = 8'd44;  #10 
a = 8'd219; b = 8'd45;  #10 
a = 8'd219; b = 8'd46;  #10 
a = 8'd219; b = 8'd47;  #10 
a = 8'd219; b = 8'd48;  #10 
a = 8'd219; b = 8'd49;  #10 
a = 8'd219; b = 8'd50;  #10 
a = 8'd219; b = 8'd51;  #10 
a = 8'd219; b = 8'd52;  #10 
a = 8'd219; b = 8'd53;  #10 
a = 8'd219; b = 8'd54;  #10 
a = 8'd219; b = 8'd55;  #10 
a = 8'd219; b = 8'd56;  #10 
a = 8'd219; b = 8'd57;  #10 
a = 8'd219; b = 8'd58;  #10 
a = 8'd219; b = 8'd59;  #10 
a = 8'd219; b = 8'd60;  #10 
a = 8'd219; b = 8'd61;  #10 
a = 8'd219; b = 8'd62;  #10 
a = 8'd219; b = 8'd63;  #10 
a = 8'd219; b = 8'd64;  #10 
a = 8'd219; b = 8'd65;  #10 
a = 8'd219; b = 8'd66;  #10 
a = 8'd219; b = 8'd67;  #10 
a = 8'd219; b = 8'd68;  #10 
a = 8'd219; b = 8'd69;  #10 
a = 8'd219; b = 8'd70;  #10 
a = 8'd219; b = 8'd71;  #10 
a = 8'd219; b = 8'd72;  #10 
a = 8'd219; b = 8'd73;  #10 
a = 8'd219; b = 8'd74;  #10 
a = 8'd219; b = 8'd75;  #10 
a = 8'd219; b = 8'd76;  #10 
a = 8'd219; b = 8'd77;  #10 
a = 8'd219; b = 8'd78;  #10 
a = 8'd219; b = 8'd79;  #10 
a = 8'd219; b = 8'd80;  #10 
a = 8'd219; b = 8'd81;  #10 
a = 8'd219; b = 8'd82;  #10 
a = 8'd219; b = 8'd83;  #10 
a = 8'd219; b = 8'd84;  #10 
a = 8'd219; b = 8'd85;  #10 
a = 8'd219; b = 8'd86;  #10 
a = 8'd219; b = 8'd87;  #10 
a = 8'd219; b = 8'd88;  #10 
a = 8'd219; b = 8'd89;  #10 
a = 8'd219; b = 8'd90;  #10 
a = 8'd219; b = 8'd91;  #10 
a = 8'd219; b = 8'd92;  #10 
a = 8'd219; b = 8'd93;  #10 
a = 8'd219; b = 8'd94;  #10 
a = 8'd219; b = 8'd95;  #10 
a = 8'd219; b = 8'd96;  #10 
a = 8'd219; b = 8'd97;  #10 
a = 8'd219; b = 8'd98;  #10 
a = 8'd219; b = 8'd99;  #10 
a = 8'd219; b = 8'd100;  #10 
a = 8'd219; b = 8'd101;  #10 
a = 8'd219; b = 8'd102;  #10 
a = 8'd219; b = 8'd103;  #10 
a = 8'd219; b = 8'd104;  #10 
a = 8'd219; b = 8'd105;  #10 
a = 8'd219; b = 8'd106;  #10 
a = 8'd219; b = 8'd107;  #10 
a = 8'd219; b = 8'd108;  #10 
a = 8'd219; b = 8'd109;  #10 
a = 8'd219; b = 8'd110;  #10 
a = 8'd219; b = 8'd111;  #10 
a = 8'd219; b = 8'd112;  #10 
a = 8'd219; b = 8'd113;  #10 
a = 8'd219; b = 8'd114;  #10 
a = 8'd219; b = 8'd115;  #10 
a = 8'd219; b = 8'd116;  #10 
a = 8'd219; b = 8'd117;  #10 
a = 8'd219; b = 8'd118;  #10 
a = 8'd219; b = 8'd119;  #10 
a = 8'd219; b = 8'd120;  #10 
a = 8'd219; b = 8'd121;  #10 
a = 8'd219; b = 8'd122;  #10 
a = 8'd219; b = 8'd123;  #10 
a = 8'd219; b = 8'd124;  #10 
a = 8'd219; b = 8'd125;  #10 
a = 8'd219; b = 8'd126;  #10 
a = 8'd219; b = 8'd127;  #10 
a = 8'd219; b = 8'd128;  #10 
a = 8'd219; b = 8'd129;  #10 
a = 8'd219; b = 8'd130;  #10 
a = 8'd219; b = 8'd131;  #10 
a = 8'd219; b = 8'd132;  #10 
a = 8'd219; b = 8'd133;  #10 
a = 8'd219; b = 8'd134;  #10 
a = 8'd219; b = 8'd135;  #10 
a = 8'd219; b = 8'd136;  #10 
a = 8'd219; b = 8'd137;  #10 
a = 8'd219; b = 8'd138;  #10 
a = 8'd219; b = 8'd139;  #10 
a = 8'd219; b = 8'd140;  #10 
a = 8'd219; b = 8'd141;  #10 
a = 8'd219; b = 8'd142;  #10 
a = 8'd219; b = 8'd143;  #10 
a = 8'd219; b = 8'd144;  #10 
a = 8'd219; b = 8'd145;  #10 
a = 8'd219; b = 8'd146;  #10 
a = 8'd219; b = 8'd147;  #10 
a = 8'd219; b = 8'd148;  #10 
a = 8'd219; b = 8'd149;  #10 
a = 8'd219; b = 8'd150;  #10 
a = 8'd219; b = 8'd151;  #10 
a = 8'd219; b = 8'd152;  #10 
a = 8'd219; b = 8'd153;  #10 
a = 8'd219; b = 8'd154;  #10 
a = 8'd219; b = 8'd155;  #10 
a = 8'd219; b = 8'd156;  #10 
a = 8'd219; b = 8'd157;  #10 
a = 8'd219; b = 8'd158;  #10 
a = 8'd219; b = 8'd159;  #10 
a = 8'd219; b = 8'd160;  #10 
a = 8'd219; b = 8'd161;  #10 
a = 8'd219; b = 8'd162;  #10 
a = 8'd219; b = 8'd163;  #10 
a = 8'd219; b = 8'd164;  #10 
a = 8'd219; b = 8'd165;  #10 
a = 8'd219; b = 8'd166;  #10 
a = 8'd219; b = 8'd167;  #10 
a = 8'd219; b = 8'd168;  #10 
a = 8'd219; b = 8'd169;  #10 
a = 8'd219; b = 8'd170;  #10 
a = 8'd219; b = 8'd171;  #10 
a = 8'd219; b = 8'd172;  #10 
a = 8'd219; b = 8'd173;  #10 
a = 8'd219; b = 8'd174;  #10 
a = 8'd219; b = 8'd175;  #10 
a = 8'd219; b = 8'd176;  #10 
a = 8'd219; b = 8'd177;  #10 
a = 8'd219; b = 8'd178;  #10 
a = 8'd219; b = 8'd179;  #10 
a = 8'd219; b = 8'd180;  #10 
a = 8'd219; b = 8'd181;  #10 
a = 8'd219; b = 8'd182;  #10 
a = 8'd219; b = 8'd183;  #10 
a = 8'd219; b = 8'd184;  #10 
a = 8'd219; b = 8'd185;  #10 
a = 8'd219; b = 8'd186;  #10 
a = 8'd219; b = 8'd187;  #10 
a = 8'd219; b = 8'd188;  #10 
a = 8'd219; b = 8'd189;  #10 
a = 8'd219; b = 8'd190;  #10 
a = 8'd219; b = 8'd191;  #10 
a = 8'd219; b = 8'd192;  #10 
a = 8'd219; b = 8'd193;  #10 
a = 8'd219; b = 8'd194;  #10 
a = 8'd219; b = 8'd195;  #10 
a = 8'd219; b = 8'd196;  #10 
a = 8'd219; b = 8'd197;  #10 
a = 8'd219; b = 8'd198;  #10 
a = 8'd219; b = 8'd199;  #10 
a = 8'd219; b = 8'd200;  #10 
a = 8'd219; b = 8'd201;  #10 
a = 8'd219; b = 8'd202;  #10 
a = 8'd219; b = 8'd203;  #10 
a = 8'd219; b = 8'd204;  #10 
a = 8'd219; b = 8'd205;  #10 
a = 8'd219; b = 8'd206;  #10 
a = 8'd219; b = 8'd207;  #10 
a = 8'd219; b = 8'd208;  #10 
a = 8'd219; b = 8'd209;  #10 
a = 8'd219; b = 8'd210;  #10 
a = 8'd219; b = 8'd211;  #10 
a = 8'd219; b = 8'd212;  #10 
a = 8'd219; b = 8'd213;  #10 
a = 8'd219; b = 8'd214;  #10 
a = 8'd219; b = 8'd215;  #10 
a = 8'd219; b = 8'd216;  #10 
a = 8'd219; b = 8'd217;  #10 
a = 8'd219; b = 8'd218;  #10 
a = 8'd219; b = 8'd219;  #10 
a = 8'd219; b = 8'd220;  #10 
a = 8'd219; b = 8'd221;  #10 
a = 8'd219; b = 8'd222;  #10 
a = 8'd219; b = 8'd223;  #10 
a = 8'd219; b = 8'd224;  #10 
a = 8'd219; b = 8'd225;  #10 
a = 8'd219; b = 8'd226;  #10 
a = 8'd219; b = 8'd227;  #10 
a = 8'd219; b = 8'd228;  #10 
a = 8'd219; b = 8'd229;  #10 
a = 8'd219; b = 8'd230;  #10 
a = 8'd219; b = 8'd231;  #10 
a = 8'd219; b = 8'd232;  #10 
a = 8'd219; b = 8'd233;  #10 
a = 8'd219; b = 8'd234;  #10 
a = 8'd219; b = 8'd235;  #10 
a = 8'd219; b = 8'd236;  #10 
a = 8'd219; b = 8'd237;  #10 
a = 8'd219; b = 8'd238;  #10 
a = 8'd219; b = 8'd239;  #10 
a = 8'd219; b = 8'd240;  #10 
a = 8'd219; b = 8'd241;  #10 
a = 8'd219; b = 8'd242;  #10 
a = 8'd219; b = 8'd243;  #10 
a = 8'd219; b = 8'd244;  #10 
a = 8'd219; b = 8'd245;  #10 
a = 8'd219; b = 8'd246;  #10 
a = 8'd219; b = 8'd247;  #10 
a = 8'd219; b = 8'd248;  #10 
a = 8'd219; b = 8'd249;  #10 
a = 8'd219; b = 8'd250;  #10 
a = 8'd219; b = 8'd251;  #10 
a = 8'd219; b = 8'd252;  #10 
a = 8'd219; b = 8'd253;  #10 
a = 8'd219; b = 8'd254;  #10 
a = 8'd219; b = 8'd255;  #10 
a = 8'd220; b = 8'd0;  #10 
a = 8'd220; b = 8'd1;  #10 
a = 8'd220; b = 8'd2;  #10 
a = 8'd220; b = 8'd3;  #10 
a = 8'd220; b = 8'd4;  #10 
a = 8'd220; b = 8'd5;  #10 
a = 8'd220; b = 8'd6;  #10 
a = 8'd220; b = 8'd7;  #10 
a = 8'd220; b = 8'd8;  #10 
a = 8'd220; b = 8'd9;  #10 
a = 8'd220; b = 8'd10;  #10 
a = 8'd220; b = 8'd11;  #10 
a = 8'd220; b = 8'd12;  #10 
a = 8'd220; b = 8'd13;  #10 
a = 8'd220; b = 8'd14;  #10 
a = 8'd220; b = 8'd15;  #10 
a = 8'd220; b = 8'd16;  #10 
a = 8'd220; b = 8'd17;  #10 
a = 8'd220; b = 8'd18;  #10 
a = 8'd220; b = 8'd19;  #10 
a = 8'd220; b = 8'd20;  #10 
a = 8'd220; b = 8'd21;  #10 
a = 8'd220; b = 8'd22;  #10 
a = 8'd220; b = 8'd23;  #10 
a = 8'd220; b = 8'd24;  #10 
a = 8'd220; b = 8'd25;  #10 
a = 8'd220; b = 8'd26;  #10 
a = 8'd220; b = 8'd27;  #10 
a = 8'd220; b = 8'd28;  #10 
a = 8'd220; b = 8'd29;  #10 
a = 8'd220; b = 8'd30;  #10 
a = 8'd220; b = 8'd31;  #10 
a = 8'd220; b = 8'd32;  #10 
a = 8'd220; b = 8'd33;  #10 
a = 8'd220; b = 8'd34;  #10 
a = 8'd220; b = 8'd35;  #10 
a = 8'd220; b = 8'd36;  #10 
a = 8'd220; b = 8'd37;  #10 
a = 8'd220; b = 8'd38;  #10 
a = 8'd220; b = 8'd39;  #10 
a = 8'd220; b = 8'd40;  #10 
a = 8'd220; b = 8'd41;  #10 
a = 8'd220; b = 8'd42;  #10 
a = 8'd220; b = 8'd43;  #10 
a = 8'd220; b = 8'd44;  #10 
a = 8'd220; b = 8'd45;  #10 
a = 8'd220; b = 8'd46;  #10 
a = 8'd220; b = 8'd47;  #10 
a = 8'd220; b = 8'd48;  #10 
a = 8'd220; b = 8'd49;  #10 
a = 8'd220; b = 8'd50;  #10 
a = 8'd220; b = 8'd51;  #10 
a = 8'd220; b = 8'd52;  #10 
a = 8'd220; b = 8'd53;  #10 
a = 8'd220; b = 8'd54;  #10 
a = 8'd220; b = 8'd55;  #10 
a = 8'd220; b = 8'd56;  #10 
a = 8'd220; b = 8'd57;  #10 
a = 8'd220; b = 8'd58;  #10 
a = 8'd220; b = 8'd59;  #10 
a = 8'd220; b = 8'd60;  #10 
a = 8'd220; b = 8'd61;  #10 
a = 8'd220; b = 8'd62;  #10 
a = 8'd220; b = 8'd63;  #10 
a = 8'd220; b = 8'd64;  #10 
a = 8'd220; b = 8'd65;  #10 
a = 8'd220; b = 8'd66;  #10 
a = 8'd220; b = 8'd67;  #10 
a = 8'd220; b = 8'd68;  #10 
a = 8'd220; b = 8'd69;  #10 
a = 8'd220; b = 8'd70;  #10 
a = 8'd220; b = 8'd71;  #10 
a = 8'd220; b = 8'd72;  #10 
a = 8'd220; b = 8'd73;  #10 
a = 8'd220; b = 8'd74;  #10 
a = 8'd220; b = 8'd75;  #10 
a = 8'd220; b = 8'd76;  #10 
a = 8'd220; b = 8'd77;  #10 
a = 8'd220; b = 8'd78;  #10 
a = 8'd220; b = 8'd79;  #10 
a = 8'd220; b = 8'd80;  #10 
a = 8'd220; b = 8'd81;  #10 
a = 8'd220; b = 8'd82;  #10 
a = 8'd220; b = 8'd83;  #10 
a = 8'd220; b = 8'd84;  #10 
a = 8'd220; b = 8'd85;  #10 
a = 8'd220; b = 8'd86;  #10 
a = 8'd220; b = 8'd87;  #10 
a = 8'd220; b = 8'd88;  #10 
a = 8'd220; b = 8'd89;  #10 
a = 8'd220; b = 8'd90;  #10 
a = 8'd220; b = 8'd91;  #10 
a = 8'd220; b = 8'd92;  #10 
a = 8'd220; b = 8'd93;  #10 
a = 8'd220; b = 8'd94;  #10 
a = 8'd220; b = 8'd95;  #10 
a = 8'd220; b = 8'd96;  #10 
a = 8'd220; b = 8'd97;  #10 
a = 8'd220; b = 8'd98;  #10 
a = 8'd220; b = 8'd99;  #10 
a = 8'd220; b = 8'd100;  #10 
a = 8'd220; b = 8'd101;  #10 
a = 8'd220; b = 8'd102;  #10 
a = 8'd220; b = 8'd103;  #10 
a = 8'd220; b = 8'd104;  #10 
a = 8'd220; b = 8'd105;  #10 
a = 8'd220; b = 8'd106;  #10 
a = 8'd220; b = 8'd107;  #10 
a = 8'd220; b = 8'd108;  #10 
a = 8'd220; b = 8'd109;  #10 
a = 8'd220; b = 8'd110;  #10 
a = 8'd220; b = 8'd111;  #10 
a = 8'd220; b = 8'd112;  #10 
a = 8'd220; b = 8'd113;  #10 
a = 8'd220; b = 8'd114;  #10 
a = 8'd220; b = 8'd115;  #10 
a = 8'd220; b = 8'd116;  #10 
a = 8'd220; b = 8'd117;  #10 
a = 8'd220; b = 8'd118;  #10 
a = 8'd220; b = 8'd119;  #10 
a = 8'd220; b = 8'd120;  #10 
a = 8'd220; b = 8'd121;  #10 
a = 8'd220; b = 8'd122;  #10 
a = 8'd220; b = 8'd123;  #10 
a = 8'd220; b = 8'd124;  #10 
a = 8'd220; b = 8'd125;  #10 
a = 8'd220; b = 8'd126;  #10 
a = 8'd220; b = 8'd127;  #10 
a = 8'd220; b = 8'd128;  #10 
a = 8'd220; b = 8'd129;  #10 
a = 8'd220; b = 8'd130;  #10 
a = 8'd220; b = 8'd131;  #10 
a = 8'd220; b = 8'd132;  #10 
a = 8'd220; b = 8'd133;  #10 
a = 8'd220; b = 8'd134;  #10 
a = 8'd220; b = 8'd135;  #10 
a = 8'd220; b = 8'd136;  #10 
a = 8'd220; b = 8'd137;  #10 
a = 8'd220; b = 8'd138;  #10 
a = 8'd220; b = 8'd139;  #10 
a = 8'd220; b = 8'd140;  #10 
a = 8'd220; b = 8'd141;  #10 
a = 8'd220; b = 8'd142;  #10 
a = 8'd220; b = 8'd143;  #10 
a = 8'd220; b = 8'd144;  #10 
a = 8'd220; b = 8'd145;  #10 
a = 8'd220; b = 8'd146;  #10 
a = 8'd220; b = 8'd147;  #10 
a = 8'd220; b = 8'd148;  #10 
a = 8'd220; b = 8'd149;  #10 
a = 8'd220; b = 8'd150;  #10 
a = 8'd220; b = 8'd151;  #10 
a = 8'd220; b = 8'd152;  #10 
a = 8'd220; b = 8'd153;  #10 
a = 8'd220; b = 8'd154;  #10 
a = 8'd220; b = 8'd155;  #10 
a = 8'd220; b = 8'd156;  #10 
a = 8'd220; b = 8'd157;  #10 
a = 8'd220; b = 8'd158;  #10 
a = 8'd220; b = 8'd159;  #10 
a = 8'd220; b = 8'd160;  #10 
a = 8'd220; b = 8'd161;  #10 
a = 8'd220; b = 8'd162;  #10 
a = 8'd220; b = 8'd163;  #10 
a = 8'd220; b = 8'd164;  #10 
a = 8'd220; b = 8'd165;  #10 
a = 8'd220; b = 8'd166;  #10 
a = 8'd220; b = 8'd167;  #10 
a = 8'd220; b = 8'd168;  #10 
a = 8'd220; b = 8'd169;  #10 
a = 8'd220; b = 8'd170;  #10 
a = 8'd220; b = 8'd171;  #10 
a = 8'd220; b = 8'd172;  #10 
a = 8'd220; b = 8'd173;  #10 
a = 8'd220; b = 8'd174;  #10 
a = 8'd220; b = 8'd175;  #10 
a = 8'd220; b = 8'd176;  #10 
a = 8'd220; b = 8'd177;  #10 
a = 8'd220; b = 8'd178;  #10 
a = 8'd220; b = 8'd179;  #10 
a = 8'd220; b = 8'd180;  #10 
a = 8'd220; b = 8'd181;  #10 
a = 8'd220; b = 8'd182;  #10 
a = 8'd220; b = 8'd183;  #10 
a = 8'd220; b = 8'd184;  #10 
a = 8'd220; b = 8'd185;  #10 
a = 8'd220; b = 8'd186;  #10 
a = 8'd220; b = 8'd187;  #10 
a = 8'd220; b = 8'd188;  #10 
a = 8'd220; b = 8'd189;  #10 
a = 8'd220; b = 8'd190;  #10 
a = 8'd220; b = 8'd191;  #10 
a = 8'd220; b = 8'd192;  #10 
a = 8'd220; b = 8'd193;  #10 
a = 8'd220; b = 8'd194;  #10 
a = 8'd220; b = 8'd195;  #10 
a = 8'd220; b = 8'd196;  #10 
a = 8'd220; b = 8'd197;  #10 
a = 8'd220; b = 8'd198;  #10 
a = 8'd220; b = 8'd199;  #10 
a = 8'd220; b = 8'd200;  #10 
a = 8'd220; b = 8'd201;  #10 
a = 8'd220; b = 8'd202;  #10 
a = 8'd220; b = 8'd203;  #10 
a = 8'd220; b = 8'd204;  #10 
a = 8'd220; b = 8'd205;  #10 
a = 8'd220; b = 8'd206;  #10 
a = 8'd220; b = 8'd207;  #10 
a = 8'd220; b = 8'd208;  #10 
a = 8'd220; b = 8'd209;  #10 
a = 8'd220; b = 8'd210;  #10 
a = 8'd220; b = 8'd211;  #10 
a = 8'd220; b = 8'd212;  #10 
a = 8'd220; b = 8'd213;  #10 
a = 8'd220; b = 8'd214;  #10 
a = 8'd220; b = 8'd215;  #10 
a = 8'd220; b = 8'd216;  #10 
a = 8'd220; b = 8'd217;  #10 
a = 8'd220; b = 8'd218;  #10 
a = 8'd220; b = 8'd219;  #10 
a = 8'd220; b = 8'd220;  #10 
a = 8'd220; b = 8'd221;  #10 
a = 8'd220; b = 8'd222;  #10 
a = 8'd220; b = 8'd223;  #10 
a = 8'd220; b = 8'd224;  #10 
a = 8'd220; b = 8'd225;  #10 
a = 8'd220; b = 8'd226;  #10 
a = 8'd220; b = 8'd227;  #10 
a = 8'd220; b = 8'd228;  #10 
a = 8'd220; b = 8'd229;  #10 
a = 8'd220; b = 8'd230;  #10 
a = 8'd220; b = 8'd231;  #10 
a = 8'd220; b = 8'd232;  #10 
a = 8'd220; b = 8'd233;  #10 
a = 8'd220; b = 8'd234;  #10 
a = 8'd220; b = 8'd235;  #10 
a = 8'd220; b = 8'd236;  #10 
a = 8'd220; b = 8'd237;  #10 
a = 8'd220; b = 8'd238;  #10 
a = 8'd220; b = 8'd239;  #10 
a = 8'd220; b = 8'd240;  #10 
a = 8'd220; b = 8'd241;  #10 
a = 8'd220; b = 8'd242;  #10 
a = 8'd220; b = 8'd243;  #10 
a = 8'd220; b = 8'd244;  #10 
a = 8'd220; b = 8'd245;  #10 
a = 8'd220; b = 8'd246;  #10 
a = 8'd220; b = 8'd247;  #10 
a = 8'd220; b = 8'd248;  #10 
a = 8'd220; b = 8'd249;  #10 
a = 8'd220; b = 8'd250;  #10 
a = 8'd220; b = 8'd251;  #10 
a = 8'd220; b = 8'd252;  #10 
a = 8'd220; b = 8'd253;  #10 
a = 8'd220; b = 8'd254;  #10 
a = 8'd220; b = 8'd255;  #10 
a = 8'd221; b = 8'd0;  #10 
a = 8'd221; b = 8'd1;  #10 
a = 8'd221; b = 8'd2;  #10 
a = 8'd221; b = 8'd3;  #10 
a = 8'd221; b = 8'd4;  #10 
a = 8'd221; b = 8'd5;  #10 
a = 8'd221; b = 8'd6;  #10 
a = 8'd221; b = 8'd7;  #10 
a = 8'd221; b = 8'd8;  #10 
a = 8'd221; b = 8'd9;  #10 
a = 8'd221; b = 8'd10;  #10 
a = 8'd221; b = 8'd11;  #10 
a = 8'd221; b = 8'd12;  #10 
a = 8'd221; b = 8'd13;  #10 
a = 8'd221; b = 8'd14;  #10 
a = 8'd221; b = 8'd15;  #10 
a = 8'd221; b = 8'd16;  #10 
a = 8'd221; b = 8'd17;  #10 
a = 8'd221; b = 8'd18;  #10 
a = 8'd221; b = 8'd19;  #10 
a = 8'd221; b = 8'd20;  #10 
a = 8'd221; b = 8'd21;  #10 
a = 8'd221; b = 8'd22;  #10 
a = 8'd221; b = 8'd23;  #10 
a = 8'd221; b = 8'd24;  #10 
a = 8'd221; b = 8'd25;  #10 
a = 8'd221; b = 8'd26;  #10 
a = 8'd221; b = 8'd27;  #10 
a = 8'd221; b = 8'd28;  #10 
a = 8'd221; b = 8'd29;  #10 
a = 8'd221; b = 8'd30;  #10 
a = 8'd221; b = 8'd31;  #10 
a = 8'd221; b = 8'd32;  #10 
a = 8'd221; b = 8'd33;  #10 
a = 8'd221; b = 8'd34;  #10 
a = 8'd221; b = 8'd35;  #10 
a = 8'd221; b = 8'd36;  #10 
a = 8'd221; b = 8'd37;  #10 
a = 8'd221; b = 8'd38;  #10 
a = 8'd221; b = 8'd39;  #10 
a = 8'd221; b = 8'd40;  #10 
a = 8'd221; b = 8'd41;  #10 
a = 8'd221; b = 8'd42;  #10 
a = 8'd221; b = 8'd43;  #10 
a = 8'd221; b = 8'd44;  #10 
a = 8'd221; b = 8'd45;  #10 
a = 8'd221; b = 8'd46;  #10 
a = 8'd221; b = 8'd47;  #10 
a = 8'd221; b = 8'd48;  #10 
a = 8'd221; b = 8'd49;  #10 
a = 8'd221; b = 8'd50;  #10 
a = 8'd221; b = 8'd51;  #10 
a = 8'd221; b = 8'd52;  #10 
a = 8'd221; b = 8'd53;  #10 
a = 8'd221; b = 8'd54;  #10 
a = 8'd221; b = 8'd55;  #10 
a = 8'd221; b = 8'd56;  #10 
a = 8'd221; b = 8'd57;  #10 
a = 8'd221; b = 8'd58;  #10 
a = 8'd221; b = 8'd59;  #10 
a = 8'd221; b = 8'd60;  #10 
a = 8'd221; b = 8'd61;  #10 
a = 8'd221; b = 8'd62;  #10 
a = 8'd221; b = 8'd63;  #10 
a = 8'd221; b = 8'd64;  #10 
a = 8'd221; b = 8'd65;  #10 
a = 8'd221; b = 8'd66;  #10 
a = 8'd221; b = 8'd67;  #10 
a = 8'd221; b = 8'd68;  #10 
a = 8'd221; b = 8'd69;  #10 
a = 8'd221; b = 8'd70;  #10 
a = 8'd221; b = 8'd71;  #10 
a = 8'd221; b = 8'd72;  #10 
a = 8'd221; b = 8'd73;  #10 
a = 8'd221; b = 8'd74;  #10 
a = 8'd221; b = 8'd75;  #10 
a = 8'd221; b = 8'd76;  #10 
a = 8'd221; b = 8'd77;  #10 
a = 8'd221; b = 8'd78;  #10 
a = 8'd221; b = 8'd79;  #10 
a = 8'd221; b = 8'd80;  #10 
a = 8'd221; b = 8'd81;  #10 
a = 8'd221; b = 8'd82;  #10 
a = 8'd221; b = 8'd83;  #10 
a = 8'd221; b = 8'd84;  #10 
a = 8'd221; b = 8'd85;  #10 
a = 8'd221; b = 8'd86;  #10 
a = 8'd221; b = 8'd87;  #10 
a = 8'd221; b = 8'd88;  #10 
a = 8'd221; b = 8'd89;  #10 
a = 8'd221; b = 8'd90;  #10 
a = 8'd221; b = 8'd91;  #10 
a = 8'd221; b = 8'd92;  #10 
a = 8'd221; b = 8'd93;  #10 
a = 8'd221; b = 8'd94;  #10 
a = 8'd221; b = 8'd95;  #10 
a = 8'd221; b = 8'd96;  #10 
a = 8'd221; b = 8'd97;  #10 
a = 8'd221; b = 8'd98;  #10 
a = 8'd221; b = 8'd99;  #10 
a = 8'd221; b = 8'd100;  #10 
a = 8'd221; b = 8'd101;  #10 
a = 8'd221; b = 8'd102;  #10 
a = 8'd221; b = 8'd103;  #10 
a = 8'd221; b = 8'd104;  #10 
a = 8'd221; b = 8'd105;  #10 
a = 8'd221; b = 8'd106;  #10 
a = 8'd221; b = 8'd107;  #10 
a = 8'd221; b = 8'd108;  #10 
a = 8'd221; b = 8'd109;  #10 
a = 8'd221; b = 8'd110;  #10 
a = 8'd221; b = 8'd111;  #10 
a = 8'd221; b = 8'd112;  #10 
a = 8'd221; b = 8'd113;  #10 
a = 8'd221; b = 8'd114;  #10 
a = 8'd221; b = 8'd115;  #10 
a = 8'd221; b = 8'd116;  #10 
a = 8'd221; b = 8'd117;  #10 
a = 8'd221; b = 8'd118;  #10 
a = 8'd221; b = 8'd119;  #10 
a = 8'd221; b = 8'd120;  #10 
a = 8'd221; b = 8'd121;  #10 
a = 8'd221; b = 8'd122;  #10 
a = 8'd221; b = 8'd123;  #10 
a = 8'd221; b = 8'd124;  #10 
a = 8'd221; b = 8'd125;  #10 
a = 8'd221; b = 8'd126;  #10 
a = 8'd221; b = 8'd127;  #10 
a = 8'd221; b = 8'd128;  #10 
a = 8'd221; b = 8'd129;  #10 
a = 8'd221; b = 8'd130;  #10 
a = 8'd221; b = 8'd131;  #10 
a = 8'd221; b = 8'd132;  #10 
a = 8'd221; b = 8'd133;  #10 
a = 8'd221; b = 8'd134;  #10 
a = 8'd221; b = 8'd135;  #10 
a = 8'd221; b = 8'd136;  #10 
a = 8'd221; b = 8'd137;  #10 
a = 8'd221; b = 8'd138;  #10 
a = 8'd221; b = 8'd139;  #10 
a = 8'd221; b = 8'd140;  #10 
a = 8'd221; b = 8'd141;  #10 
a = 8'd221; b = 8'd142;  #10 
a = 8'd221; b = 8'd143;  #10 
a = 8'd221; b = 8'd144;  #10 
a = 8'd221; b = 8'd145;  #10 
a = 8'd221; b = 8'd146;  #10 
a = 8'd221; b = 8'd147;  #10 
a = 8'd221; b = 8'd148;  #10 
a = 8'd221; b = 8'd149;  #10 
a = 8'd221; b = 8'd150;  #10 
a = 8'd221; b = 8'd151;  #10 
a = 8'd221; b = 8'd152;  #10 
a = 8'd221; b = 8'd153;  #10 
a = 8'd221; b = 8'd154;  #10 
a = 8'd221; b = 8'd155;  #10 
a = 8'd221; b = 8'd156;  #10 
a = 8'd221; b = 8'd157;  #10 
a = 8'd221; b = 8'd158;  #10 
a = 8'd221; b = 8'd159;  #10 
a = 8'd221; b = 8'd160;  #10 
a = 8'd221; b = 8'd161;  #10 
a = 8'd221; b = 8'd162;  #10 
a = 8'd221; b = 8'd163;  #10 
a = 8'd221; b = 8'd164;  #10 
a = 8'd221; b = 8'd165;  #10 
a = 8'd221; b = 8'd166;  #10 
a = 8'd221; b = 8'd167;  #10 
a = 8'd221; b = 8'd168;  #10 
a = 8'd221; b = 8'd169;  #10 
a = 8'd221; b = 8'd170;  #10 
a = 8'd221; b = 8'd171;  #10 
a = 8'd221; b = 8'd172;  #10 
a = 8'd221; b = 8'd173;  #10 
a = 8'd221; b = 8'd174;  #10 
a = 8'd221; b = 8'd175;  #10 
a = 8'd221; b = 8'd176;  #10 
a = 8'd221; b = 8'd177;  #10 
a = 8'd221; b = 8'd178;  #10 
a = 8'd221; b = 8'd179;  #10 
a = 8'd221; b = 8'd180;  #10 
a = 8'd221; b = 8'd181;  #10 
a = 8'd221; b = 8'd182;  #10 
a = 8'd221; b = 8'd183;  #10 
a = 8'd221; b = 8'd184;  #10 
a = 8'd221; b = 8'd185;  #10 
a = 8'd221; b = 8'd186;  #10 
a = 8'd221; b = 8'd187;  #10 
a = 8'd221; b = 8'd188;  #10 
a = 8'd221; b = 8'd189;  #10 
a = 8'd221; b = 8'd190;  #10 
a = 8'd221; b = 8'd191;  #10 
a = 8'd221; b = 8'd192;  #10 
a = 8'd221; b = 8'd193;  #10 
a = 8'd221; b = 8'd194;  #10 
a = 8'd221; b = 8'd195;  #10 
a = 8'd221; b = 8'd196;  #10 
a = 8'd221; b = 8'd197;  #10 
a = 8'd221; b = 8'd198;  #10 
a = 8'd221; b = 8'd199;  #10 
a = 8'd221; b = 8'd200;  #10 
a = 8'd221; b = 8'd201;  #10 
a = 8'd221; b = 8'd202;  #10 
a = 8'd221; b = 8'd203;  #10 
a = 8'd221; b = 8'd204;  #10 
a = 8'd221; b = 8'd205;  #10 
a = 8'd221; b = 8'd206;  #10 
a = 8'd221; b = 8'd207;  #10 
a = 8'd221; b = 8'd208;  #10 
a = 8'd221; b = 8'd209;  #10 
a = 8'd221; b = 8'd210;  #10 
a = 8'd221; b = 8'd211;  #10 
a = 8'd221; b = 8'd212;  #10 
a = 8'd221; b = 8'd213;  #10 
a = 8'd221; b = 8'd214;  #10 
a = 8'd221; b = 8'd215;  #10 
a = 8'd221; b = 8'd216;  #10 
a = 8'd221; b = 8'd217;  #10 
a = 8'd221; b = 8'd218;  #10 
a = 8'd221; b = 8'd219;  #10 
a = 8'd221; b = 8'd220;  #10 
a = 8'd221; b = 8'd221;  #10 
a = 8'd221; b = 8'd222;  #10 
a = 8'd221; b = 8'd223;  #10 
a = 8'd221; b = 8'd224;  #10 
a = 8'd221; b = 8'd225;  #10 
a = 8'd221; b = 8'd226;  #10 
a = 8'd221; b = 8'd227;  #10 
a = 8'd221; b = 8'd228;  #10 
a = 8'd221; b = 8'd229;  #10 
a = 8'd221; b = 8'd230;  #10 
a = 8'd221; b = 8'd231;  #10 
a = 8'd221; b = 8'd232;  #10 
a = 8'd221; b = 8'd233;  #10 
a = 8'd221; b = 8'd234;  #10 
a = 8'd221; b = 8'd235;  #10 
a = 8'd221; b = 8'd236;  #10 
a = 8'd221; b = 8'd237;  #10 
a = 8'd221; b = 8'd238;  #10 
a = 8'd221; b = 8'd239;  #10 
a = 8'd221; b = 8'd240;  #10 
a = 8'd221; b = 8'd241;  #10 
a = 8'd221; b = 8'd242;  #10 
a = 8'd221; b = 8'd243;  #10 
a = 8'd221; b = 8'd244;  #10 
a = 8'd221; b = 8'd245;  #10 
a = 8'd221; b = 8'd246;  #10 
a = 8'd221; b = 8'd247;  #10 
a = 8'd221; b = 8'd248;  #10 
a = 8'd221; b = 8'd249;  #10 
a = 8'd221; b = 8'd250;  #10 
a = 8'd221; b = 8'd251;  #10 
a = 8'd221; b = 8'd252;  #10 
a = 8'd221; b = 8'd253;  #10 
a = 8'd221; b = 8'd254;  #10 
a = 8'd221; b = 8'd255;  #10 
a = 8'd222; b = 8'd0;  #10 
a = 8'd222; b = 8'd1;  #10 
a = 8'd222; b = 8'd2;  #10 
a = 8'd222; b = 8'd3;  #10 
a = 8'd222; b = 8'd4;  #10 
a = 8'd222; b = 8'd5;  #10 
a = 8'd222; b = 8'd6;  #10 
a = 8'd222; b = 8'd7;  #10 
a = 8'd222; b = 8'd8;  #10 
a = 8'd222; b = 8'd9;  #10 
a = 8'd222; b = 8'd10;  #10 
a = 8'd222; b = 8'd11;  #10 
a = 8'd222; b = 8'd12;  #10 
a = 8'd222; b = 8'd13;  #10 
a = 8'd222; b = 8'd14;  #10 
a = 8'd222; b = 8'd15;  #10 
a = 8'd222; b = 8'd16;  #10 
a = 8'd222; b = 8'd17;  #10 
a = 8'd222; b = 8'd18;  #10 
a = 8'd222; b = 8'd19;  #10 
a = 8'd222; b = 8'd20;  #10 
a = 8'd222; b = 8'd21;  #10 
a = 8'd222; b = 8'd22;  #10 
a = 8'd222; b = 8'd23;  #10 
a = 8'd222; b = 8'd24;  #10 
a = 8'd222; b = 8'd25;  #10 
a = 8'd222; b = 8'd26;  #10 
a = 8'd222; b = 8'd27;  #10 
a = 8'd222; b = 8'd28;  #10 
a = 8'd222; b = 8'd29;  #10 
a = 8'd222; b = 8'd30;  #10 
a = 8'd222; b = 8'd31;  #10 
a = 8'd222; b = 8'd32;  #10 
a = 8'd222; b = 8'd33;  #10 
a = 8'd222; b = 8'd34;  #10 
a = 8'd222; b = 8'd35;  #10 
a = 8'd222; b = 8'd36;  #10 
a = 8'd222; b = 8'd37;  #10 
a = 8'd222; b = 8'd38;  #10 
a = 8'd222; b = 8'd39;  #10 
a = 8'd222; b = 8'd40;  #10 
a = 8'd222; b = 8'd41;  #10 
a = 8'd222; b = 8'd42;  #10 
a = 8'd222; b = 8'd43;  #10 
a = 8'd222; b = 8'd44;  #10 
a = 8'd222; b = 8'd45;  #10 
a = 8'd222; b = 8'd46;  #10 
a = 8'd222; b = 8'd47;  #10 
a = 8'd222; b = 8'd48;  #10 
a = 8'd222; b = 8'd49;  #10 
a = 8'd222; b = 8'd50;  #10 
a = 8'd222; b = 8'd51;  #10 
a = 8'd222; b = 8'd52;  #10 
a = 8'd222; b = 8'd53;  #10 
a = 8'd222; b = 8'd54;  #10 
a = 8'd222; b = 8'd55;  #10 
a = 8'd222; b = 8'd56;  #10 
a = 8'd222; b = 8'd57;  #10 
a = 8'd222; b = 8'd58;  #10 
a = 8'd222; b = 8'd59;  #10 
a = 8'd222; b = 8'd60;  #10 
a = 8'd222; b = 8'd61;  #10 
a = 8'd222; b = 8'd62;  #10 
a = 8'd222; b = 8'd63;  #10 
a = 8'd222; b = 8'd64;  #10 
a = 8'd222; b = 8'd65;  #10 
a = 8'd222; b = 8'd66;  #10 
a = 8'd222; b = 8'd67;  #10 
a = 8'd222; b = 8'd68;  #10 
a = 8'd222; b = 8'd69;  #10 
a = 8'd222; b = 8'd70;  #10 
a = 8'd222; b = 8'd71;  #10 
a = 8'd222; b = 8'd72;  #10 
a = 8'd222; b = 8'd73;  #10 
a = 8'd222; b = 8'd74;  #10 
a = 8'd222; b = 8'd75;  #10 
a = 8'd222; b = 8'd76;  #10 
a = 8'd222; b = 8'd77;  #10 
a = 8'd222; b = 8'd78;  #10 
a = 8'd222; b = 8'd79;  #10 
a = 8'd222; b = 8'd80;  #10 
a = 8'd222; b = 8'd81;  #10 
a = 8'd222; b = 8'd82;  #10 
a = 8'd222; b = 8'd83;  #10 
a = 8'd222; b = 8'd84;  #10 
a = 8'd222; b = 8'd85;  #10 
a = 8'd222; b = 8'd86;  #10 
a = 8'd222; b = 8'd87;  #10 
a = 8'd222; b = 8'd88;  #10 
a = 8'd222; b = 8'd89;  #10 
a = 8'd222; b = 8'd90;  #10 
a = 8'd222; b = 8'd91;  #10 
a = 8'd222; b = 8'd92;  #10 
a = 8'd222; b = 8'd93;  #10 
a = 8'd222; b = 8'd94;  #10 
a = 8'd222; b = 8'd95;  #10 
a = 8'd222; b = 8'd96;  #10 
a = 8'd222; b = 8'd97;  #10 
a = 8'd222; b = 8'd98;  #10 
a = 8'd222; b = 8'd99;  #10 
a = 8'd222; b = 8'd100;  #10 
a = 8'd222; b = 8'd101;  #10 
a = 8'd222; b = 8'd102;  #10 
a = 8'd222; b = 8'd103;  #10 
a = 8'd222; b = 8'd104;  #10 
a = 8'd222; b = 8'd105;  #10 
a = 8'd222; b = 8'd106;  #10 
a = 8'd222; b = 8'd107;  #10 
a = 8'd222; b = 8'd108;  #10 
a = 8'd222; b = 8'd109;  #10 
a = 8'd222; b = 8'd110;  #10 
a = 8'd222; b = 8'd111;  #10 
a = 8'd222; b = 8'd112;  #10 
a = 8'd222; b = 8'd113;  #10 
a = 8'd222; b = 8'd114;  #10 
a = 8'd222; b = 8'd115;  #10 
a = 8'd222; b = 8'd116;  #10 
a = 8'd222; b = 8'd117;  #10 
a = 8'd222; b = 8'd118;  #10 
a = 8'd222; b = 8'd119;  #10 
a = 8'd222; b = 8'd120;  #10 
a = 8'd222; b = 8'd121;  #10 
a = 8'd222; b = 8'd122;  #10 
a = 8'd222; b = 8'd123;  #10 
a = 8'd222; b = 8'd124;  #10 
a = 8'd222; b = 8'd125;  #10 
a = 8'd222; b = 8'd126;  #10 
a = 8'd222; b = 8'd127;  #10 
a = 8'd222; b = 8'd128;  #10 
a = 8'd222; b = 8'd129;  #10 
a = 8'd222; b = 8'd130;  #10 
a = 8'd222; b = 8'd131;  #10 
a = 8'd222; b = 8'd132;  #10 
a = 8'd222; b = 8'd133;  #10 
a = 8'd222; b = 8'd134;  #10 
a = 8'd222; b = 8'd135;  #10 
a = 8'd222; b = 8'd136;  #10 
a = 8'd222; b = 8'd137;  #10 
a = 8'd222; b = 8'd138;  #10 
a = 8'd222; b = 8'd139;  #10 
a = 8'd222; b = 8'd140;  #10 
a = 8'd222; b = 8'd141;  #10 
a = 8'd222; b = 8'd142;  #10 
a = 8'd222; b = 8'd143;  #10 
a = 8'd222; b = 8'd144;  #10 
a = 8'd222; b = 8'd145;  #10 
a = 8'd222; b = 8'd146;  #10 
a = 8'd222; b = 8'd147;  #10 
a = 8'd222; b = 8'd148;  #10 
a = 8'd222; b = 8'd149;  #10 
a = 8'd222; b = 8'd150;  #10 
a = 8'd222; b = 8'd151;  #10 
a = 8'd222; b = 8'd152;  #10 
a = 8'd222; b = 8'd153;  #10 
a = 8'd222; b = 8'd154;  #10 
a = 8'd222; b = 8'd155;  #10 
a = 8'd222; b = 8'd156;  #10 
a = 8'd222; b = 8'd157;  #10 
a = 8'd222; b = 8'd158;  #10 
a = 8'd222; b = 8'd159;  #10 
a = 8'd222; b = 8'd160;  #10 
a = 8'd222; b = 8'd161;  #10 
a = 8'd222; b = 8'd162;  #10 
a = 8'd222; b = 8'd163;  #10 
a = 8'd222; b = 8'd164;  #10 
a = 8'd222; b = 8'd165;  #10 
a = 8'd222; b = 8'd166;  #10 
a = 8'd222; b = 8'd167;  #10 
a = 8'd222; b = 8'd168;  #10 
a = 8'd222; b = 8'd169;  #10 
a = 8'd222; b = 8'd170;  #10 
a = 8'd222; b = 8'd171;  #10 
a = 8'd222; b = 8'd172;  #10 
a = 8'd222; b = 8'd173;  #10 
a = 8'd222; b = 8'd174;  #10 
a = 8'd222; b = 8'd175;  #10 
a = 8'd222; b = 8'd176;  #10 
a = 8'd222; b = 8'd177;  #10 
a = 8'd222; b = 8'd178;  #10 
a = 8'd222; b = 8'd179;  #10 
a = 8'd222; b = 8'd180;  #10 
a = 8'd222; b = 8'd181;  #10 
a = 8'd222; b = 8'd182;  #10 
a = 8'd222; b = 8'd183;  #10 
a = 8'd222; b = 8'd184;  #10 
a = 8'd222; b = 8'd185;  #10 
a = 8'd222; b = 8'd186;  #10 
a = 8'd222; b = 8'd187;  #10 
a = 8'd222; b = 8'd188;  #10 
a = 8'd222; b = 8'd189;  #10 
a = 8'd222; b = 8'd190;  #10 
a = 8'd222; b = 8'd191;  #10 
a = 8'd222; b = 8'd192;  #10 
a = 8'd222; b = 8'd193;  #10 
a = 8'd222; b = 8'd194;  #10 
a = 8'd222; b = 8'd195;  #10 
a = 8'd222; b = 8'd196;  #10 
a = 8'd222; b = 8'd197;  #10 
a = 8'd222; b = 8'd198;  #10 
a = 8'd222; b = 8'd199;  #10 
a = 8'd222; b = 8'd200;  #10 
a = 8'd222; b = 8'd201;  #10 
a = 8'd222; b = 8'd202;  #10 
a = 8'd222; b = 8'd203;  #10 
a = 8'd222; b = 8'd204;  #10 
a = 8'd222; b = 8'd205;  #10 
a = 8'd222; b = 8'd206;  #10 
a = 8'd222; b = 8'd207;  #10 
a = 8'd222; b = 8'd208;  #10 
a = 8'd222; b = 8'd209;  #10 
a = 8'd222; b = 8'd210;  #10 
a = 8'd222; b = 8'd211;  #10 
a = 8'd222; b = 8'd212;  #10 
a = 8'd222; b = 8'd213;  #10 
a = 8'd222; b = 8'd214;  #10 
a = 8'd222; b = 8'd215;  #10 
a = 8'd222; b = 8'd216;  #10 
a = 8'd222; b = 8'd217;  #10 
a = 8'd222; b = 8'd218;  #10 
a = 8'd222; b = 8'd219;  #10 
a = 8'd222; b = 8'd220;  #10 
a = 8'd222; b = 8'd221;  #10 
a = 8'd222; b = 8'd222;  #10 
a = 8'd222; b = 8'd223;  #10 
a = 8'd222; b = 8'd224;  #10 
a = 8'd222; b = 8'd225;  #10 
a = 8'd222; b = 8'd226;  #10 
a = 8'd222; b = 8'd227;  #10 
a = 8'd222; b = 8'd228;  #10 
a = 8'd222; b = 8'd229;  #10 
a = 8'd222; b = 8'd230;  #10 
a = 8'd222; b = 8'd231;  #10 
a = 8'd222; b = 8'd232;  #10 
a = 8'd222; b = 8'd233;  #10 
a = 8'd222; b = 8'd234;  #10 
a = 8'd222; b = 8'd235;  #10 
a = 8'd222; b = 8'd236;  #10 
a = 8'd222; b = 8'd237;  #10 
a = 8'd222; b = 8'd238;  #10 
a = 8'd222; b = 8'd239;  #10 
a = 8'd222; b = 8'd240;  #10 
a = 8'd222; b = 8'd241;  #10 
a = 8'd222; b = 8'd242;  #10 
a = 8'd222; b = 8'd243;  #10 
a = 8'd222; b = 8'd244;  #10 
a = 8'd222; b = 8'd245;  #10 
a = 8'd222; b = 8'd246;  #10 
a = 8'd222; b = 8'd247;  #10 
a = 8'd222; b = 8'd248;  #10 
a = 8'd222; b = 8'd249;  #10 
a = 8'd222; b = 8'd250;  #10 
a = 8'd222; b = 8'd251;  #10 
a = 8'd222; b = 8'd252;  #10 
a = 8'd222; b = 8'd253;  #10 
a = 8'd222; b = 8'd254;  #10 
a = 8'd222; b = 8'd255;  #10 
a = 8'd223; b = 8'd0;  #10 
a = 8'd223; b = 8'd1;  #10 
a = 8'd223; b = 8'd2;  #10 
a = 8'd223; b = 8'd3;  #10 
a = 8'd223; b = 8'd4;  #10 
a = 8'd223; b = 8'd5;  #10 
a = 8'd223; b = 8'd6;  #10 
a = 8'd223; b = 8'd7;  #10 
a = 8'd223; b = 8'd8;  #10 
a = 8'd223; b = 8'd9;  #10 
a = 8'd223; b = 8'd10;  #10 
a = 8'd223; b = 8'd11;  #10 
a = 8'd223; b = 8'd12;  #10 
a = 8'd223; b = 8'd13;  #10 
a = 8'd223; b = 8'd14;  #10 
a = 8'd223; b = 8'd15;  #10 
a = 8'd223; b = 8'd16;  #10 
a = 8'd223; b = 8'd17;  #10 
a = 8'd223; b = 8'd18;  #10 
a = 8'd223; b = 8'd19;  #10 
a = 8'd223; b = 8'd20;  #10 
a = 8'd223; b = 8'd21;  #10 
a = 8'd223; b = 8'd22;  #10 
a = 8'd223; b = 8'd23;  #10 
a = 8'd223; b = 8'd24;  #10 
a = 8'd223; b = 8'd25;  #10 
a = 8'd223; b = 8'd26;  #10 
a = 8'd223; b = 8'd27;  #10 
a = 8'd223; b = 8'd28;  #10 
a = 8'd223; b = 8'd29;  #10 
a = 8'd223; b = 8'd30;  #10 
a = 8'd223; b = 8'd31;  #10 
a = 8'd223; b = 8'd32;  #10 
a = 8'd223; b = 8'd33;  #10 
a = 8'd223; b = 8'd34;  #10 
a = 8'd223; b = 8'd35;  #10 
a = 8'd223; b = 8'd36;  #10 
a = 8'd223; b = 8'd37;  #10 
a = 8'd223; b = 8'd38;  #10 
a = 8'd223; b = 8'd39;  #10 
a = 8'd223; b = 8'd40;  #10 
a = 8'd223; b = 8'd41;  #10 
a = 8'd223; b = 8'd42;  #10 
a = 8'd223; b = 8'd43;  #10 
a = 8'd223; b = 8'd44;  #10 
a = 8'd223; b = 8'd45;  #10 
a = 8'd223; b = 8'd46;  #10 
a = 8'd223; b = 8'd47;  #10 
a = 8'd223; b = 8'd48;  #10 
a = 8'd223; b = 8'd49;  #10 
a = 8'd223; b = 8'd50;  #10 
a = 8'd223; b = 8'd51;  #10 
a = 8'd223; b = 8'd52;  #10 
a = 8'd223; b = 8'd53;  #10 
a = 8'd223; b = 8'd54;  #10 
a = 8'd223; b = 8'd55;  #10 
a = 8'd223; b = 8'd56;  #10 
a = 8'd223; b = 8'd57;  #10 
a = 8'd223; b = 8'd58;  #10 
a = 8'd223; b = 8'd59;  #10 
a = 8'd223; b = 8'd60;  #10 
a = 8'd223; b = 8'd61;  #10 
a = 8'd223; b = 8'd62;  #10 
a = 8'd223; b = 8'd63;  #10 
a = 8'd223; b = 8'd64;  #10 
a = 8'd223; b = 8'd65;  #10 
a = 8'd223; b = 8'd66;  #10 
a = 8'd223; b = 8'd67;  #10 
a = 8'd223; b = 8'd68;  #10 
a = 8'd223; b = 8'd69;  #10 
a = 8'd223; b = 8'd70;  #10 
a = 8'd223; b = 8'd71;  #10 
a = 8'd223; b = 8'd72;  #10 
a = 8'd223; b = 8'd73;  #10 
a = 8'd223; b = 8'd74;  #10 
a = 8'd223; b = 8'd75;  #10 
a = 8'd223; b = 8'd76;  #10 
a = 8'd223; b = 8'd77;  #10 
a = 8'd223; b = 8'd78;  #10 
a = 8'd223; b = 8'd79;  #10 
a = 8'd223; b = 8'd80;  #10 
a = 8'd223; b = 8'd81;  #10 
a = 8'd223; b = 8'd82;  #10 
a = 8'd223; b = 8'd83;  #10 
a = 8'd223; b = 8'd84;  #10 
a = 8'd223; b = 8'd85;  #10 
a = 8'd223; b = 8'd86;  #10 
a = 8'd223; b = 8'd87;  #10 
a = 8'd223; b = 8'd88;  #10 
a = 8'd223; b = 8'd89;  #10 
a = 8'd223; b = 8'd90;  #10 
a = 8'd223; b = 8'd91;  #10 
a = 8'd223; b = 8'd92;  #10 
a = 8'd223; b = 8'd93;  #10 
a = 8'd223; b = 8'd94;  #10 
a = 8'd223; b = 8'd95;  #10 
a = 8'd223; b = 8'd96;  #10 
a = 8'd223; b = 8'd97;  #10 
a = 8'd223; b = 8'd98;  #10 
a = 8'd223; b = 8'd99;  #10 
a = 8'd223; b = 8'd100;  #10 
a = 8'd223; b = 8'd101;  #10 
a = 8'd223; b = 8'd102;  #10 
a = 8'd223; b = 8'd103;  #10 
a = 8'd223; b = 8'd104;  #10 
a = 8'd223; b = 8'd105;  #10 
a = 8'd223; b = 8'd106;  #10 
a = 8'd223; b = 8'd107;  #10 
a = 8'd223; b = 8'd108;  #10 
a = 8'd223; b = 8'd109;  #10 
a = 8'd223; b = 8'd110;  #10 
a = 8'd223; b = 8'd111;  #10 
a = 8'd223; b = 8'd112;  #10 
a = 8'd223; b = 8'd113;  #10 
a = 8'd223; b = 8'd114;  #10 
a = 8'd223; b = 8'd115;  #10 
a = 8'd223; b = 8'd116;  #10 
a = 8'd223; b = 8'd117;  #10 
a = 8'd223; b = 8'd118;  #10 
a = 8'd223; b = 8'd119;  #10 
a = 8'd223; b = 8'd120;  #10 
a = 8'd223; b = 8'd121;  #10 
a = 8'd223; b = 8'd122;  #10 
a = 8'd223; b = 8'd123;  #10 
a = 8'd223; b = 8'd124;  #10 
a = 8'd223; b = 8'd125;  #10 
a = 8'd223; b = 8'd126;  #10 
a = 8'd223; b = 8'd127;  #10 
a = 8'd223; b = 8'd128;  #10 
a = 8'd223; b = 8'd129;  #10 
a = 8'd223; b = 8'd130;  #10 
a = 8'd223; b = 8'd131;  #10 
a = 8'd223; b = 8'd132;  #10 
a = 8'd223; b = 8'd133;  #10 
a = 8'd223; b = 8'd134;  #10 
a = 8'd223; b = 8'd135;  #10 
a = 8'd223; b = 8'd136;  #10 
a = 8'd223; b = 8'd137;  #10 
a = 8'd223; b = 8'd138;  #10 
a = 8'd223; b = 8'd139;  #10 
a = 8'd223; b = 8'd140;  #10 
a = 8'd223; b = 8'd141;  #10 
a = 8'd223; b = 8'd142;  #10 
a = 8'd223; b = 8'd143;  #10 
a = 8'd223; b = 8'd144;  #10 
a = 8'd223; b = 8'd145;  #10 
a = 8'd223; b = 8'd146;  #10 
a = 8'd223; b = 8'd147;  #10 
a = 8'd223; b = 8'd148;  #10 
a = 8'd223; b = 8'd149;  #10 
a = 8'd223; b = 8'd150;  #10 
a = 8'd223; b = 8'd151;  #10 
a = 8'd223; b = 8'd152;  #10 
a = 8'd223; b = 8'd153;  #10 
a = 8'd223; b = 8'd154;  #10 
a = 8'd223; b = 8'd155;  #10 
a = 8'd223; b = 8'd156;  #10 
a = 8'd223; b = 8'd157;  #10 
a = 8'd223; b = 8'd158;  #10 
a = 8'd223; b = 8'd159;  #10 
a = 8'd223; b = 8'd160;  #10 
a = 8'd223; b = 8'd161;  #10 
a = 8'd223; b = 8'd162;  #10 
a = 8'd223; b = 8'd163;  #10 
a = 8'd223; b = 8'd164;  #10 
a = 8'd223; b = 8'd165;  #10 
a = 8'd223; b = 8'd166;  #10 
a = 8'd223; b = 8'd167;  #10 
a = 8'd223; b = 8'd168;  #10 
a = 8'd223; b = 8'd169;  #10 
a = 8'd223; b = 8'd170;  #10 
a = 8'd223; b = 8'd171;  #10 
a = 8'd223; b = 8'd172;  #10 
a = 8'd223; b = 8'd173;  #10 
a = 8'd223; b = 8'd174;  #10 
a = 8'd223; b = 8'd175;  #10 
a = 8'd223; b = 8'd176;  #10 
a = 8'd223; b = 8'd177;  #10 
a = 8'd223; b = 8'd178;  #10 
a = 8'd223; b = 8'd179;  #10 
a = 8'd223; b = 8'd180;  #10 
a = 8'd223; b = 8'd181;  #10 
a = 8'd223; b = 8'd182;  #10 
a = 8'd223; b = 8'd183;  #10 
a = 8'd223; b = 8'd184;  #10 
a = 8'd223; b = 8'd185;  #10 
a = 8'd223; b = 8'd186;  #10 
a = 8'd223; b = 8'd187;  #10 
a = 8'd223; b = 8'd188;  #10 
a = 8'd223; b = 8'd189;  #10 
a = 8'd223; b = 8'd190;  #10 
a = 8'd223; b = 8'd191;  #10 
a = 8'd223; b = 8'd192;  #10 
a = 8'd223; b = 8'd193;  #10 
a = 8'd223; b = 8'd194;  #10 
a = 8'd223; b = 8'd195;  #10 
a = 8'd223; b = 8'd196;  #10 
a = 8'd223; b = 8'd197;  #10 
a = 8'd223; b = 8'd198;  #10 
a = 8'd223; b = 8'd199;  #10 
a = 8'd223; b = 8'd200;  #10 
a = 8'd223; b = 8'd201;  #10 
a = 8'd223; b = 8'd202;  #10 
a = 8'd223; b = 8'd203;  #10 
a = 8'd223; b = 8'd204;  #10 
a = 8'd223; b = 8'd205;  #10 
a = 8'd223; b = 8'd206;  #10 
a = 8'd223; b = 8'd207;  #10 
a = 8'd223; b = 8'd208;  #10 
a = 8'd223; b = 8'd209;  #10 
a = 8'd223; b = 8'd210;  #10 
a = 8'd223; b = 8'd211;  #10 
a = 8'd223; b = 8'd212;  #10 
a = 8'd223; b = 8'd213;  #10 
a = 8'd223; b = 8'd214;  #10 
a = 8'd223; b = 8'd215;  #10 
a = 8'd223; b = 8'd216;  #10 
a = 8'd223; b = 8'd217;  #10 
a = 8'd223; b = 8'd218;  #10 
a = 8'd223; b = 8'd219;  #10 
a = 8'd223; b = 8'd220;  #10 
a = 8'd223; b = 8'd221;  #10 
a = 8'd223; b = 8'd222;  #10 
a = 8'd223; b = 8'd223;  #10 
a = 8'd223; b = 8'd224;  #10 
a = 8'd223; b = 8'd225;  #10 
a = 8'd223; b = 8'd226;  #10 
a = 8'd223; b = 8'd227;  #10 
a = 8'd223; b = 8'd228;  #10 
a = 8'd223; b = 8'd229;  #10 
a = 8'd223; b = 8'd230;  #10 
a = 8'd223; b = 8'd231;  #10 
a = 8'd223; b = 8'd232;  #10 
a = 8'd223; b = 8'd233;  #10 
a = 8'd223; b = 8'd234;  #10 
a = 8'd223; b = 8'd235;  #10 
a = 8'd223; b = 8'd236;  #10 
a = 8'd223; b = 8'd237;  #10 
a = 8'd223; b = 8'd238;  #10 
a = 8'd223; b = 8'd239;  #10 
a = 8'd223; b = 8'd240;  #10 
a = 8'd223; b = 8'd241;  #10 
a = 8'd223; b = 8'd242;  #10 
a = 8'd223; b = 8'd243;  #10 
a = 8'd223; b = 8'd244;  #10 
a = 8'd223; b = 8'd245;  #10 
a = 8'd223; b = 8'd246;  #10 
a = 8'd223; b = 8'd247;  #10 
a = 8'd223; b = 8'd248;  #10 
a = 8'd223; b = 8'd249;  #10 
a = 8'd223; b = 8'd250;  #10 
a = 8'd223; b = 8'd251;  #10 
a = 8'd223; b = 8'd252;  #10 
a = 8'd223; b = 8'd253;  #10 
a = 8'd223; b = 8'd254;  #10 
a = 8'd223; b = 8'd255;  #10 
a = 8'd224; b = 8'd0;  #10 
a = 8'd224; b = 8'd1;  #10 
a = 8'd224; b = 8'd2;  #10 
a = 8'd224; b = 8'd3;  #10 
a = 8'd224; b = 8'd4;  #10 
a = 8'd224; b = 8'd5;  #10 
a = 8'd224; b = 8'd6;  #10 
a = 8'd224; b = 8'd7;  #10 
a = 8'd224; b = 8'd8;  #10 
a = 8'd224; b = 8'd9;  #10 
a = 8'd224; b = 8'd10;  #10 
a = 8'd224; b = 8'd11;  #10 
a = 8'd224; b = 8'd12;  #10 
a = 8'd224; b = 8'd13;  #10 
a = 8'd224; b = 8'd14;  #10 
a = 8'd224; b = 8'd15;  #10 
a = 8'd224; b = 8'd16;  #10 
a = 8'd224; b = 8'd17;  #10 
a = 8'd224; b = 8'd18;  #10 
a = 8'd224; b = 8'd19;  #10 
a = 8'd224; b = 8'd20;  #10 
a = 8'd224; b = 8'd21;  #10 
a = 8'd224; b = 8'd22;  #10 
a = 8'd224; b = 8'd23;  #10 
a = 8'd224; b = 8'd24;  #10 
a = 8'd224; b = 8'd25;  #10 
a = 8'd224; b = 8'd26;  #10 
a = 8'd224; b = 8'd27;  #10 
a = 8'd224; b = 8'd28;  #10 
a = 8'd224; b = 8'd29;  #10 
a = 8'd224; b = 8'd30;  #10 
a = 8'd224; b = 8'd31;  #10 
a = 8'd224; b = 8'd32;  #10 
a = 8'd224; b = 8'd33;  #10 
a = 8'd224; b = 8'd34;  #10 
a = 8'd224; b = 8'd35;  #10 
a = 8'd224; b = 8'd36;  #10 
a = 8'd224; b = 8'd37;  #10 
a = 8'd224; b = 8'd38;  #10 
a = 8'd224; b = 8'd39;  #10 
a = 8'd224; b = 8'd40;  #10 
a = 8'd224; b = 8'd41;  #10 
a = 8'd224; b = 8'd42;  #10 
a = 8'd224; b = 8'd43;  #10 
a = 8'd224; b = 8'd44;  #10 
a = 8'd224; b = 8'd45;  #10 
a = 8'd224; b = 8'd46;  #10 
a = 8'd224; b = 8'd47;  #10 
a = 8'd224; b = 8'd48;  #10 
a = 8'd224; b = 8'd49;  #10 
a = 8'd224; b = 8'd50;  #10 
a = 8'd224; b = 8'd51;  #10 
a = 8'd224; b = 8'd52;  #10 
a = 8'd224; b = 8'd53;  #10 
a = 8'd224; b = 8'd54;  #10 
a = 8'd224; b = 8'd55;  #10 
a = 8'd224; b = 8'd56;  #10 
a = 8'd224; b = 8'd57;  #10 
a = 8'd224; b = 8'd58;  #10 
a = 8'd224; b = 8'd59;  #10 
a = 8'd224; b = 8'd60;  #10 
a = 8'd224; b = 8'd61;  #10 
a = 8'd224; b = 8'd62;  #10 
a = 8'd224; b = 8'd63;  #10 
a = 8'd224; b = 8'd64;  #10 
a = 8'd224; b = 8'd65;  #10 
a = 8'd224; b = 8'd66;  #10 
a = 8'd224; b = 8'd67;  #10 
a = 8'd224; b = 8'd68;  #10 
a = 8'd224; b = 8'd69;  #10 
a = 8'd224; b = 8'd70;  #10 
a = 8'd224; b = 8'd71;  #10 
a = 8'd224; b = 8'd72;  #10 
a = 8'd224; b = 8'd73;  #10 
a = 8'd224; b = 8'd74;  #10 
a = 8'd224; b = 8'd75;  #10 
a = 8'd224; b = 8'd76;  #10 
a = 8'd224; b = 8'd77;  #10 
a = 8'd224; b = 8'd78;  #10 
a = 8'd224; b = 8'd79;  #10 
a = 8'd224; b = 8'd80;  #10 
a = 8'd224; b = 8'd81;  #10 
a = 8'd224; b = 8'd82;  #10 
a = 8'd224; b = 8'd83;  #10 
a = 8'd224; b = 8'd84;  #10 
a = 8'd224; b = 8'd85;  #10 
a = 8'd224; b = 8'd86;  #10 
a = 8'd224; b = 8'd87;  #10 
a = 8'd224; b = 8'd88;  #10 
a = 8'd224; b = 8'd89;  #10 
a = 8'd224; b = 8'd90;  #10 
a = 8'd224; b = 8'd91;  #10 
a = 8'd224; b = 8'd92;  #10 
a = 8'd224; b = 8'd93;  #10 
a = 8'd224; b = 8'd94;  #10 
a = 8'd224; b = 8'd95;  #10 
a = 8'd224; b = 8'd96;  #10 
a = 8'd224; b = 8'd97;  #10 
a = 8'd224; b = 8'd98;  #10 
a = 8'd224; b = 8'd99;  #10 
a = 8'd224; b = 8'd100;  #10 
a = 8'd224; b = 8'd101;  #10 
a = 8'd224; b = 8'd102;  #10 
a = 8'd224; b = 8'd103;  #10 
a = 8'd224; b = 8'd104;  #10 
a = 8'd224; b = 8'd105;  #10 
a = 8'd224; b = 8'd106;  #10 
a = 8'd224; b = 8'd107;  #10 
a = 8'd224; b = 8'd108;  #10 
a = 8'd224; b = 8'd109;  #10 
a = 8'd224; b = 8'd110;  #10 
a = 8'd224; b = 8'd111;  #10 
a = 8'd224; b = 8'd112;  #10 
a = 8'd224; b = 8'd113;  #10 
a = 8'd224; b = 8'd114;  #10 
a = 8'd224; b = 8'd115;  #10 
a = 8'd224; b = 8'd116;  #10 
a = 8'd224; b = 8'd117;  #10 
a = 8'd224; b = 8'd118;  #10 
a = 8'd224; b = 8'd119;  #10 
a = 8'd224; b = 8'd120;  #10 
a = 8'd224; b = 8'd121;  #10 
a = 8'd224; b = 8'd122;  #10 
a = 8'd224; b = 8'd123;  #10 
a = 8'd224; b = 8'd124;  #10 
a = 8'd224; b = 8'd125;  #10 
a = 8'd224; b = 8'd126;  #10 
a = 8'd224; b = 8'd127;  #10 
a = 8'd224; b = 8'd128;  #10 
a = 8'd224; b = 8'd129;  #10 
a = 8'd224; b = 8'd130;  #10 
a = 8'd224; b = 8'd131;  #10 
a = 8'd224; b = 8'd132;  #10 
a = 8'd224; b = 8'd133;  #10 
a = 8'd224; b = 8'd134;  #10 
a = 8'd224; b = 8'd135;  #10 
a = 8'd224; b = 8'd136;  #10 
a = 8'd224; b = 8'd137;  #10 
a = 8'd224; b = 8'd138;  #10 
a = 8'd224; b = 8'd139;  #10 
a = 8'd224; b = 8'd140;  #10 
a = 8'd224; b = 8'd141;  #10 
a = 8'd224; b = 8'd142;  #10 
a = 8'd224; b = 8'd143;  #10 
a = 8'd224; b = 8'd144;  #10 
a = 8'd224; b = 8'd145;  #10 
a = 8'd224; b = 8'd146;  #10 
a = 8'd224; b = 8'd147;  #10 
a = 8'd224; b = 8'd148;  #10 
a = 8'd224; b = 8'd149;  #10 
a = 8'd224; b = 8'd150;  #10 
a = 8'd224; b = 8'd151;  #10 
a = 8'd224; b = 8'd152;  #10 
a = 8'd224; b = 8'd153;  #10 
a = 8'd224; b = 8'd154;  #10 
a = 8'd224; b = 8'd155;  #10 
a = 8'd224; b = 8'd156;  #10 
a = 8'd224; b = 8'd157;  #10 
a = 8'd224; b = 8'd158;  #10 
a = 8'd224; b = 8'd159;  #10 
a = 8'd224; b = 8'd160;  #10 
a = 8'd224; b = 8'd161;  #10 
a = 8'd224; b = 8'd162;  #10 
a = 8'd224; b = 8'd163;  #10 
a = 8'd224; b = 8'd164;  #10 
a = 8'd224; b = 8'd165;  #10 
a = 8'd224; b = 8'd166;  #10 
a = 8'd224; b = 8'd167;  #10 
a = 8'd224; b = 8'd168;  #10 
a = 8'd224; b = 8'd169;  #10 
a = 8'd224; b = 8'd170;  #10 
a = 8'd224; b = 8'd171;  #10 
a = 8'd224; b = 8'd172;  #10 
a = 8'd224; b = 8'd173;  #10 
a = 8'd224; b = 8'd174;  #10 
a = 8'd224; b = 8'd175;  #10 
a = 8'd224; b = 8'd176;  #10 
a = 8'd224; b = 8'd177;  #10 
a = 8'd224; b = 8'd178;  #10 
a = 8'd224; b = 8'd179;  #10 
a = 8'd224; b = 8'd180;  #10 
a = 8'd224; b = 8'd181;  #10 
a = 8'd224; b = 8'd182;  #10 
a = 8'd224; b = 8'd183;  #10 
a = 8'd224; b = 8'd184;  #10 
a = 8'd224; b = 8'd185;  #10 
a = 8'd224; b = 8'd186;  #10 
a = 8'd224; b = 8'd187;  #10 
a = 8'd224; b = 8'd188;  #10 
a = 8'd224; b = 8'd189;  #10 
a = 8'd224; b = 8'd190;  #10 
a = 8'd224; b = 8'd191;  #10 
a = 8'd224; b = 8'd192;  #10 
a = 8'd224; b = 8'd193;  #10 
a = 8'd224; b = 8'd194;  #10 
a = 8'd224; b = 8'd195;  #10 
a = 8'd224; b = 8'd196;  #10 
a = 8'd224; b = 8'd197;  #10 
a = 8'd224; b = 8'd198;  #10 
a = 8'd224; b = 8'd199;  #10 
a = 8'd224; b = 8'd200;  #10 
a = 8'd224; b = 8'd201;  #10 
a = 8'd224; b = 8'd202;  #10 
a = 8'd224; b = 8'd203;  #10 
a = 8'd224; b = 8'd204;  #10 
a = 8'd224; b = 8'd205;  #10 
a = 8'd224; b = 8'd206;  #10 
a = 8'd224; b = 8'd207;  #10 
a = 8'd224; b = 8'd208;  #10 
a = 8'd224; b = 8'd209;  #10 
a = 8'd224; b = 8'd210;  #10 
a = 8'd224; b = 8'd211;  #10 
a = 8'd224; b = 8'd212;  #10 
a = 8'd224; b = 8'd213;  #10 
a = 8'd224; b = 8'd214;  #10 
a = 8'd224; b = 8'd215;  #10 
a = 8'd224; b = 8'd216;  #10 
a = 8'd224; b = 8'd217;  #10 
a = 8'd224; b = 8'd218;  #10 
a = 8'd224; b = 8'd219;  #10 
a = 8'd224; b = 8'd220;  #10 
a = 8'd224; b = 8'd221;  #10 
a = 8'd224; b = 8'd222;  #10 
a = 8'd224; b = 8'd223;  #10 
a = 8'd224; b = 8'd224;  #10 
a = 8'd224; b = 8'd225;  #10 
a = 8'd224; b = 8'd226;  #10 
a = 8'd224; b = 8'd227;  #10 
a = 8'd224; b = 8'd228;  #10 
a = 8'd224; b = 8'd229;  #10 
a = 8'd224; b = 8'd230;  #10 
a = 8'd224; b = 8'd231;  #10 
a = 8'd224; b = 8'd232;  #10 
a = 8'd224; b = 8'd233;  #10 
a = 8'd224; b = 8'd234;  #10 
a = 8'd224; b = 8'd235;  #10 
a = 8'd224; b = 8'd236;  #10 
a = 8'd224; b = 8'd237;  #10 
a = 8'd224; b = 8'd238;  #10 
a = 8'd224; b = 8'd239;  #10 
a = 8'd224; b = 8'd240;  #10 
a = 8'd224; b = 8'd241;  #10 
a = 8'd224; b = 8'd242;  #10 
a = 8'd224; b = 8'd243;  #10 
a = 8'd224; b = 8'd244;  #10 
a = 8'd224; b = 8'd245;  #10 
a = 8'd224; b = 8'd246;  #10 
a = 8'd224; b = 8'd247;  #10 
a = 8'd224; b = 8'd248;  #10 
a = 8'd224; b = 8'd249;  #10 
a = 8'd224; b = 8'd250;  #10 
a = 8'd224; b = 8'd251;  #10 
a = 8'd224; b = 8'd252;  #10 
a = 8'd224; b = 8'd253;  #10 
a = 8'd224; b = 8'd254;  #10 
a = 8'd224; b = 8'd255;  #10 
a = 8'd225; b = 8'd0;  #10 
a = 8'd225; b = 8'd1;  #10 
a = 8'd225; b = 8'd2;  #10 
a = 8'd225; b = 8'd3;  #10 
a = 8'd225; b = 8'd4;  #10 
a = 8'd225; b = 8'd5;  #10 
a = 8'd225; b = 8'd6;  #10 
a = 8'd225; b = 8'd7;  #10 
a = 8'd225; b = 8'd8;  #10 
a = 8'd225; b = 8'd9;  #10 
a = 8'd225; b = 8'd10;  #10 
a = 8'd225; b = 8'd11;  #10 
a = 8'd225; b = 8'd12;  #10 
a = 8'd225; b = 8'd13;  #10 
a = 8'd225; b = 8'd14;  #10 
a = 8'd225; b = 8'd15;  #10 
a = 8'd225; b = 8'd16;  #10 
a = 8'd225; b = 8'd17;  #10 
a = 8'd225; b = 8'd18;  #10 
a = 8'd225; b = 8'd19;  #10 
a = 8'd225; b = 8'd20;  #10 
a = 8'd225; b = 8'd21;  #10 
a = 8'd225; b = 8'd22;  #10 
a = 8'd225; b = 8'd23;  #10 
a = 8'd225; b = 8'd24;  #10 
a = 8'd225; b = 8'd25;  #10 
a = 8'd225; b = 8'd26;  #10 
a = 8'd225; b = 8'd27;  #10 
a = 8'd225; b = 8'd28;  #10 
a = 8'd225; b = 8'd29;  #10 
a = 8'd225; b = 8'd30;  #10 
a = 8'd225; b = 8'd31;  #10 
a = 8'd225; b = 8'd32;  #10 
a = 8'd225; b = 8'd33;  #10 
a = 8'd225; b = 8'd34;  #10 
a = 8'd225; b = 8'd35;  #10 
a = 8'd225; b = 8'd36;  #10 
a = 8'd225; b = 8'd37;  #10 
a = 8'd225; b = 8'd38;  #10 
a = 8'd225; b = 8'd39;  #10 
a = 8'd225; b = 8'd40;  #10 
a = 8'd225; b = 8'd41;  #10 
a = 8'd225; b = 8'd42;  #10 
a = 8'd225; b = 8'd43;  #10 
a = 8'd225; b = 8'd44;  #10 
a = 8'd225; b = 8'd45;  #10 
a = 8'd225; b = 8'd46;  #10 
a = 8'd225; b = 8'd47;  #10 
a = 8'd225; b = 8'd48;  #10 
a = 8'd225; b = 8'd49;  #10 
a = 8'd225; b = 8'd50;  #10 
a = 8'd225; b = 8'd51;  #10 
a = 8'd225; b = 8'd52;  #10 
a = 8'd225; b = 8'd53;  #10 
a = 8'd225; b = 8'd54;  #10 
a = 8'd225; b = 8'd55;  #10 
a = 8'd225; b = 8'd56;  #10 
a = 8'd225; b = 8'd57;  #10 
a = 8'd225; b = 8'd58;  #10 
a = 8'd225; b = 8'd59;  #10 
a = 8'd225; b = 8'd60;  #10 
a = 8'd225; b = 8'd61;  #10 
a = 8'd225; b = 8'd62;  #10 
a = 8'd225; b = 8'd63;  #10 
a = 8'd225; b = 8'd64;  #10 
a = 8'd225; b = 8'd65;  #10 
a = 8'd225; b = 8'd66;  #10 
a = 8'd225; b = 8'd67;  #10 
a = 8'd225; b = 8'd68;  #10 
a = 8'd225; b = 8'd69;  #10 
a = 8'd225; b = 8'd70;  #10 
a = 8'd225; b = 8'd71;  #10 
a = 8'd225; b = 8'd72;  #10 
a = 8'd225; b = 8'd73;  #10 
a = 8'd225; b = 8'd74;  #10 
a = 8'd225; b = 8'd75;  #10 
a = 8'd225; b = 8'd76;  #10 
a = 8'd225; b = 8'd77;  #10 
a = 8'd225; b = 8'd78;  #10 
a = 8'd225; b = 8'd79;  #10 
a = 8'd225; b = 8'd80;  #10 
a = 8'd225; b = 8'd81;  #10 
a = 8'd225; b = 8'd82;  #10 
a = 8'd225; b = 8'd83;  #10 
a = 8'd225; b = 8'd84;  #10 
a = 8'd225; b = 8'd85;  #10 
a = 8'd225; b = 8'd86;  #10 
a = 8'd225; b = 8'd87;  #10 
a = 8'd225; b = 8'd88;  #10 
a = 8'd225; b = 8'd89;  #10 
a = 8'd225; b = 8'd90;  #10 
a = 8'd225; b = 8'd91;  #10 
a = 8'd225; b = 8'd92;  #10 
a = 8'd225; b = 8'd93;  #10 
a = 8'd225; b = 8'd94;  #10 
a = 8'd225; b = 8'd95;  #10 
a = 8'd225; b = 8'd96;  #10 
a = 8'd225; b = 8'd97;  #10 
a = 8'd225; b = 8'd98;  #10 
a = 8'd225; b = 8'd99;  #10 
a = 8'd225; b = 8'd100;  #10 
a = 8'd225; b = 8'd101;  #10 
a = 8'd225; b = 8'd102;  #10 
a = 8'd225; b = 8'd103;  #10 
a = 8'd225; b = 8'd104;  #10 
a = 8'd225; b = 8'd105;  #10 
a = 8'd225; b = 8'd106;  #10 
a = 8'd225; b = 8'd107;  #10 
a = 8'd225; b = 8'd108;  #10 
a = 8'd225; b = 8'd109;  #10 
a = 8'd225; b = 8'd110;  #10 
a = 8'd225; b = 8'd111;  #10 
a = 8'd225; b = 8'd112;  #10 
a = 8'd225; b = 8'd113;  #10 
a = 8'd225; b = 8'd114;  #10 
a = 8'd225; b = 8'd115;  #10 
a = 8'd225; b = 8'd116;  #10 
a = 8'd225; b = 8'd117;  #10 
a = 8'd225; b = 8'd118;  #10 
a = 8'd225; b = 8'd119;  #10 
a = 8'd225; b = 8'd120;  #10 
a = 8'd225; b = 8'd121;  #10 
a = 8'd225; b = 8'd122;  #10 
a = 8'd225; b = 8'd123;  #10 
a = 8'd225; b = 8'd124;  #10 
a = 8'd225; b = 8'd125;  #10 
a = 8'd225; b = 8'd126;  #10 
a = 8'd225; b = 8'd127;  #10 
a = 8'd225; b = 8'd128;  #10 
a = 8'd225; b = 8'd129;  #10 
a = 8'd225; b = 8'd130;  #10 
a = 8'd225; b = 8'd131;  #10 
a = 8'd225; b = 8'd132;  #10 
a = 8'd225; b = 8'd133;  #10 
a = 8'd225; b = 8'd134;  #10 
a = 8'd225; b = 8'd135;  #10 
a = 8'd225; b = 8'd136;  #10 
a = 8'd225; b = 8'd137;  #10 
a = 8'd225; b = 8'd138;  #10 
a = 8'd225; b = 8'd139;  #10 
a = 8'd225; b = 8'd140;  #10 
a = 8'd225; b = 8'd141;  #10 
a = 8'd225; b = 8'd142;  #10 
a = 8'd225; b = 8'd143;  #10 
a = 8'd225; b = 8'd144;  #10 
a = 8'd225; b = 8'd145;  #10 
a = 8'd225; b = 8'd146;  #10 
a = 8'd225; b = 8'd147;  #10 
a = 8'd225; b = 8'd148;  #10 
a = 8'd225; b = 8'd149;  #10 
a = 8'd225; b = 8'd150;  #10 
a = 8'd225; b = 8'd151;  #10 
a = 8'd225; b = 8'd152;  #10 
a = 8'd225; b = 8'd153;  #10 
a = 8'd225; b = 8'd154;  #10 
a = 8'd225; b = 8'd155;  #10 
a = 8'd225; b = 8'd156;  #10 
a = 8'd225; b = 8'd157;  #10 
a = 8'd225; b = 8'd158;  #10 
a = 8'd225; b = 8'd159;  #10 
a = 8'd225; b = 8'd160;  #10 
a = 8'd225; b = 8'd161;  #10 
a = 8'd225; b = 8'd162;  #10 
a = 8'd225; b = 8'd163;  #10 
a = 8'd225; b = 8'd164;  #10 
a = 8'd225; b = 8'd165;  #10 
a = 8'd225; b = 8'd166;  #10 
a = 8'd225; b = 8'd167;  #10 
a = 8'd225; b = 8'd168;  #10 
a = 8'd225; b = 8'd169;  #10 
a = 8'd225; b = 8'd170;  #10 
a = 8'd225; b = 8'd171;  #10 
a = 8'd225; b = 8'd172;  #10 
a = 8'd225; b = 8'd173;  #10 
a = 8'd225; b = 8'd174;  #10 
a = 8'd225; b = 8'd175;  #10 
a = 8'd225; b = 8'd176;  #10 
a = 8'd225; b = 8'd177;  #10 
a = 8'd225; b = 8'd178;  #10 
a = 8'd225; b = 8'd179;  #10 
a = 8'd225; b = 8'd180;  #10 
a = 8'd225; b = 8'd181;  #10 
a = 8'd225; b = 8'd182;  #10 
a = 8'd225; b = 8'd183;  #10 
a = 8'd225; b = 8'd184;  #10 
a = 8'd225; b = 8'd185;  #10 
a = 8'd225; b = 8'd186;  #10 
a = 8'd225; b = 8'd187;  #10 
a = 8'd225; b = 8'd188;  #10 
a = 8'd225; b = 8'd189;  #10 
a = 8'd225; b = 8'd190;  #10 
a = 8'd225; b = 8'd191;  #10 
a = 8'd225; b = 8'd192;  #10 
a = 8'd225; b = 8'd193;  #10 
a = 8'd225; b = 8'd194;  #10 
a = 8'd225; b = 8'd195;  #10 
a = 8'd225; b = 8'd196;  #10 
a = 8'd225; b = 8'd197;  #10 
a = 8'd225; b = 8'd198;  #10 
a = 8'd225; b = 8'd199;  #10 
a = 8'd225; b = 8'd200;  #10 
a = 8'd225; b = 8'd201;  #10 
a = 8'd225; b = 8'd202;  #10 
a = 8'd225; b = 8'd203;  #10 
a = 8'd225; b = 8'd204;  #10 
a = 8'd225; b = 8'd205;  #10 
a = 8'd225; b = 8'd206;  #10 
a = 8'd225; b = 8'd207;  #10 
a = 8'd225; b = 8'd208;  #10 
a = 8'd225; b = 8'd209;  #10 
a = 8'd225; b = 8'd210;  #10 
a = 8'd225; b = 8'd211;  #10 
a = 8'd225; b = 8'd212;  #10 
a = 8'd225; b = 8'd213;  #10 
a = 8'd225; b = 8'd214;  #10 
a = 8'd225; b = 8'd215;  #10 
a = 8'd225; b = 8'd216;  #10 
a = 8'd225; b = 8'd217;  #10 
a = 8'd225; b = 8'd218;  #10 
a = 8'd225; b = 8'd219;  #10 
a = 8'd225; b = 8'd220;  #10 
a = 8'd225; b = 8'd221;  #10 
a = 8'd225; b = 8'd222;  #10 
a = 8'd225; b = 8'd223;  #10 
a = 8'd225; b = 8'd224;  #10 
a = 8'd225; b = 8'd225;  #10 
a = 8'd225; b = 8'd226;  #10 
a = 8'd225; b = 8'd227;  #10 
a = 8'd225; b = 8'd228;  #10 
a = 8'd225; b = 8'd229;  #10 
a = 8'd225; b = 8'd230;  #10 
a = 8'd225; b = 8'd231;  #10 
a = 8'd225; b = 8'd232;  #10 
a = 8'd225; b = 8'd233;  #10 
a = 8'd225; b = 8'd234;  #10 
a = 8'd225; b = 8'd235;  #10 
a = 8'd225; b = 8'd236;  #10 
a = 8'd225; b = 8'd237;  #10 
a = 8'd225; b = 8'd238;  #10 
a = 8'd225; b = 8'd239;  #10 
a = 8'd225; b = 8'd240;  #10 
a = 8'd225; b = 8'd241;  #10 
a = 8'd225; b = 8'd242;  #10 
a = 8'd225; b = 8'd243;  #10 
a = 8'd225; b = 8'd244;  #10 
a = 8'd225; b = 8'd245;  #10 
a = 8'd225; b = 8'd246;  #10 
a = 8'd225; b = 8'd247;  #10 
a = 8'd225; b = 8'd248;  #10 
a = 8'd225; b = 8'd249;  #10 
a = 8'd225; b = 8'd250;  #10 
a = 8'd225; b = 8'd251;  #10 
a = 8'd225; b = 8'd252;  #10 
a = 8'd225; b = 8'd253;  #10 
a = 8'd225; b = 8'd254;  #10 
a = 8'd225; b = 8'd255;  #10 
a = 8'd226; b = 8'd0;  #10 
a = 8'd226; b = 8'd1;  #10 
a = 8'd226; b = 8'd2;  #10 
a = 8'd226; b = 8'd3;  #10 
a = 8'd226; b = 8'd4;  #10 
a = 8'd226; b = 8'd5;  #10 
a = 8'd226; b = 8'd6;  #10 
a = 8'd226; b = 8'd7;  #10 
a = 8'd226; b = 8'd8;  #10 
a = 8'd226; b = 8'd9;  #10 
a = 8'd226; b = 8'd10;  #10 
a = 8'd226; b = 8'd11;  #10 
a = 8'd226; b = 8'd12;  #10 
a = 8'd226; b = 8'd13;  #10 
a = 8'd226; b = 8'd14;  #10 
a = 8'd226; b = 8'd15;  #10 
a = 8'd226; b = 8'd16;  #10 
a = 8'd226; b = 8'd17;  #10 
a = 8'd226; b = 8'd18;  #10 
a = 8'd226; b = 8'd19;  #10 
a = 8'd226; b = 8'd20;  #10 
a = 8'd226; b = 8'd21;  #10 
a = 8'd226; b = 8'd22;  #10 
a = 8'd226; b = 8'd23;  #10 
a = 8'd226; b = 8'd24;  #10 
a = 8'd226; b = 8'd25;  #10 
a = 8'd226; b = 8'd26;  #10 
a = 8'd226; b = 8'd27;  #10 
a = 8'd226; b = 8'd28;  #10 
a = 8'd226; b = 8'd29;  #10 
a = 8'd226; b = 8'd30;  #10 
a = 8'd226; b = 8'd31;  #10 
a = 8'd226; b = 8'd32;  #10 
a = 8'd226; b = 8'd33;  #10 
a = 8'd226; b = 8'd34;  #10 
a = 8'd226; b = 8'd35;  #10 
a = 8'd226; b = 8'd36;  #10 
a = 8'd226; b = 8'd37;  #10 
a = 8'd226; b = 8'd38;  #10 
a = 8'd226; b = 8'd39;  #10 
a = 8'd226; b = 8'd40;  #10 
a = 8'd226; b = 8'd41;  #10 
a = 8'd226; b = 8'd42;  #10 
a = 8'd226; b = 8'd43;  #10 
a = 8'd226; b = 8'd44;  #10 
a = 8'd226; b = 8'd45;  #10 
a = 8'd226; b = 8'd46;  #10 
a = 8'd226; b = 8'd47;  #10 
a = 8'd226; b = 8'd48;  #10 
a = 8'd226; b = 8'd49;  #10 
a = 8'd226; b = 8'd50;  #10 
a = 8'd226; b = 8'd51;  #10 
a = 8'd226; b = 8'd52;  #10 
a = 8'd226; b = 8'd53;  #10 
a = 8'd226; b = 8'd54;  #10 
a = 8'd226; b = 8'd55;  #10 
a = 8'd226; b = 8'd56;  #10 
a = 8'd226; b = 8'd57;  #10 
a = 8'd226; b = 8'd58;  #10 
a = 8'd226; b = 8'd59;  #10 
a = 8'd226; b = 8'd60;  #10 
a = 8'd226; b = 8'd61;  #10 
a = 8'd226; b = 8'd62;  #10 
a = 8'd226; b = 8'd63;  #10 
a = 8'd226; b = 8'd64;  #10 
a = 8'd226; b = 8'd65;  #10 
a = 8'd226; b = 8'd66;  #10 
a = 8'd226; b = 8'd67;  #10 
a = 8'd226; b = 8'd68;  #10 
a = 8'd226; b = 8'd69;  #10 
a = 8'd226; b = 8'd70;  #10 
a = 8'd226; b = 8'd71;  #10 
a = 8'd226; b = 8'd72;  #10 
a = 8'd226; b = 8'd73;  #10 
a = 8'd226; b = 8'd74;  #10 
a = 8'd226; b = 8'd75;  #10 
a = 8'd226; b = 8'd76;  #10 
a = 8'd226; b = 8'd77;  #10 
a = 8'd226; b = 8'd78;  #10 
a = 8'd226; b = 8'd79;  #10 
a = 8'd226; b = 8'd80;  #10 
a = 8'd226; b = 8'd81;  #10 
a = 8'd226; b = 8'd82;  #10 
a = 8'd226; b = 8'd83;  #10 
a = 8'd226; b = 8'd84;  #10 
a = 8'd226; b = 8'd85;  #10 
a = 8'd226; b = 8'd86;  #10 
a = 8'd226; b = 8'd87;  #10 
a = 8'd226; b = 8'd88;  #10 
a = 8'd226; b = 8'd89;  #10 
a = 8'd226; b = 8'd90;  #10 
a = 8'd226; b = 8'd91;  #10 
a = 8'd226; b = 8'd92;  #10 
a = 8'd226; b = 8'd93;  #10 
a = 8'd226; b = 8'd94;  #10 
a = 8'd226; b = 8'd95;  #10 
a = 8'd226; b = 8'd96;  #10 
a = 8'd226; b = 8'd97;  #10 
a = 8'd226; b = 8'd98;  #10 
a = 8'd226; b = 8'd99;  #10 
a = 8'd226; b = 8'd100;  #10 
a = 8'd226; b = 8'd101;  #10 
a = 8'd226; b = 8'd102;  #10 
a = 8'd226; b = 8'd103;  #10 
a = 8'd226; b = 8'd104;  #10 
a = 8'd226; b = 8'd105;  #10 
a = 8'd226; b = 8'd106;  #10 
a = 8'd226; b = 8'd107;  #10 
a = 8'd226; b = 8'd108;  #10 
a = 8'd226; b = 8'd109;  #10 
a = 8'd226; b = 8'd110;  #10 
a = 8'd226; b = 8'd111;  #10 
a = 8'd226; b = 8'd112;  #10 
a = 8'd226; b = 8'd113;  #10 
a = 8'd226; b = 8'd114;  #10 
a = 8'd226; b = 8'd115;  #10 
a = 8'd226; b = 8'd116;  #10 
a = 8'd226; b = 8'd117;  #10 
a = 8'd226; b = 8'd118;  #10 
a = 8'd226; b = 8'd119;  #10 
a = 8'd226; b = 8'd120;  #10 
a = 8'd226; b = 8'd121;  #10 
a = 8'd226; b = 8'd122;  #10 
a = 8'd226; b = 8'd123;  #10 
a = 8'd226; b = 8'd124;  #10 
a = 8'd226; b = 8'd125;  #10 
a = 8'd226; b = 8'd126;  #10 
a = 8'd226; b = 8'd127;  #10 
a = 8'd226; b = 8'd128;  #10 
a = 8'd226; b = 8'd129;  #10 
a = 8'd226; b = 8'd130;  #10 
a = 8'd226; b = 8'd131;  #10 
a = 8'd226; b = 8'd132;  #10 
a = 8'd226; b = 8'd133;  #10 
a = 8'd226; b = 8'd134;  #10 
a = 8'd226; b = 8'd135;  #10 
a = 8'd226; b = 8'd136;  #10 
a = 8'd226; b = 8'd137;  #10 
a = 8'd226; b = 8'd138;  #10 
a = 8'd226; b = 8'd139;  #10 
a = 8'd226; b = 8'd140;  #10 
a = 8'd226; b = 8'd141;  #10 
a = 8'd226; b = 8'd142;  #10 
a = 8'd226; b = 8'd143;  #10 
a = 8'd226; b = 8'd144;  #10 
a = 8'd226; b = 8'd145;  #10 
a = 8'd226; b = 8'd146;  #10 
a = 8'd226; b = 8'd147;  #10 
a = 8'd226; b = 8'd148;  #10 
a = 8'd226; b = 8'd149;  #10 
a = 8'd226; b = 8'd150;  #10 
a = 8'd226; b = 8'd151;  #10 
a = 8'd226; b = 8'd152;  #10 
a = 8'd226; b = 8'd153;  #10 
a = 8'd226; b = 8'd154;  #10 
a = 8'd226; b = 8'd155;  #10 
a = 8'd226; b = 8'd156;  #10 
a = 8'd226; b = 8'd157;  #10 
a = 8'd226; b = 8'd158;  #10 
a = 8'd226; b = 8'd159;  #10 
a = 8'd226; b = 8'd160;  #10 
a = 8'd226; b = 8'd161;  #10 
a = 8'd226; b = 8'd162;  #10 
a = 8'd226; b = 8'd163;  #10 
a = 8'd226; b = 8'd164;  #10 
a = 8'd226; b = 8'd165;  #10 
a = 8'd226; b = 8'd166;  #10 
a = 8'd226; b = 8'd167;  #10 
a = 8'd226; b = 8'd168;  #10 
a = 8'd226; b = 8'd169;  #10 
a = 8'd226; b = 8'd170;  #10 
a = 8'd226; b = 8'd171;  #10 
a = 8'd226; b = 8'd172;  #10 
a = 8'd226; b = 8'd173;  #10 
a = 8'd226; b = 8'd174;  #10 
a = 8'd226; b = 8'd175;  #10 
a = 8'd226; b = 8'd176;  #10 
a = 8'd226; b = 8'd177;  #10 
a = 8'd226; b = 8'd178;  #10 
a = 8'd226; b = 8'd179;  #10 
a = 8'd226; b = 8'd180;  #10 
a = 8'd226; b = 8'd181;  #10 
a = 8'd226; b = 8'd182;  #10 
a = 8'd226; b = 8'd183;  #10 
a = 8'd226; b = 8'd184;  #10 
a = 8'd226; b = 8'd185;  #10 
a = 8'd226; b = 8'd186;  #10 
a = 8'd226; b = 8'd187;  #10 
a = 8'd226; b = 8'd188;  #10 
a = 8'd226; b = 8'd189;  #10 
a = 8'd226; b = 8'd190;  #10 
a = 8'd226; b = 8'd191;  #10 
a = 8'd226; b = 8'd192;  #10 
a = 8'd226; b = 8'd193;  #10 
a = 8'd226; b = 8'd194;  #10 
a = 8'd226; b = 8'd195;  #10 
a = 8'd226; b = 8'd196;  #10 
a = 8'd226; b = 8'd197;  #10 
a = 8'd226; b = 8'd198;  #10 
a = 8'd226; b = 8'd199;  #10 
a = 8'd226; b = 8'd200;  #10 
a = 8'd226; b = 8'd201;  #10 
a = 8'd226; b = 8'd202;  #10 
a = 8'd226; b = 8'd203;  #10 
a = 8'd226; b = 8'd204;  #10 
a = 8'd226; b = 8'd205;  #10 
a = 8'd226; b = 8'd206;  #10 
a = 8'd226; b = 8'd207;  #10 
a = 8'd226; b = 8'd208;  #10 
a = 8'd226; b = 8'd209;  #10 
a = 8'd226; b = 8'd210;  #10 
a = 8'd226; b = 8'd211;  #10 
a = 8'd226; b = 8'd212;  #10 
a = 8'd226; b = 8'd213;  #10 
a = 8'd226; b = 8'd214;  #10 
a = 8'd226; b = 8'd215;  #10 
a = 8'd226; b = 8'd216;  #10 
a = 8'd226; b = 8'd217;  #10 
a = 8'd226; b = 8'd218;  #10 
a = 8'd226; b = 8'd219;  #10 
a = 8'd226; b = 8'd220;  #10 
a = 8'd226; b = 8'd221;  #10 
a = 8'd226; b = 8'd222;  #10 
a = 8'd226; b = 8'd223;  #10 
a = 8'd226; b = 8'd224;  #10 
a = 8'd226; b = 8'd225;  #10 
a = 8'd226; b = 8'd226;  #10 
a = 8'd226; b = 8'd227;  #10 
a = 8'd226; b = 8'd228;  #10 
a = 8'd226; b = 8'd229;  #10 
a = 8'd226; b = 8'd230;  #10 
a = 8'd226; b = 8'd231;  #10 
a = 8'd226; b = 8'd232;  #10 
a = 8'd226; b = 8'd233;  #10 
a = 8'd226; b = 8'd234;  #10 
a = 8'd226; b = 8'd235;  #10 
a = 8'd226; b = 8'd236;  #10 
a = 8'd226; b = 8'd237;  #10 
a = 8'd226; b = 8'd238;  #10 
a = 8'd226; b = 8'd239;  #10 
a = 8'd226; b = 8'd240;  #10 
a = 8'd226; b = 8'd241;  #10 
a = 8'd226; b = 8'd242;  #10 
a = 8'd226; b = 8'd243;  #10 
a = 8'd226; b = 8'd244;  #10 
a = 8'd226; b = 8'd245;  #10 
a = 8'd226; b = 8'd246;  #10 
a = 8'd226; b = 8'd247;  #10 
a = 8'd226; b = 8'd248;  #10 
a = 8'd226; b = 8'd249;  #10 
a = 8'd226; b = 8'd250;  #10 
a = 8'd226; b = 8'd251;  #10 
a = 8'd226; b = 8'd252;  #10 
a = 8'd226; b = 8'd253;  #10 
a = 8'd226; b = 8'd254;  #10 
a = 8'd226; b = 8'd255;  #10 
a = 8'd227; b = 8'd0;  #10 
a = 8'd227; b = 8'd1;  #10 
a = 8'd227; b = 8'd2;  #10 
a = 8'd227; b = 8'd3;  #10 
a = 8'd227; b = 8'd4;  #10 
a = 8'd227; b = 8'd5;  #10 
a = 8'd227; b = 8'd6;  #10 
a = 8'd227; b = 8'd7;  #10 
a = 8'd227; b = 8'd8;  #10 
a = 8'd227; b = 8'd9;  #10 
a = 8'd227; b = 8'd10;  #10 
a = 8'd227; b = 8'd11;  #10 
a = 8'd227; b = 8'd12;  #10 
a = 8'd227; b = 8'd13;  #10 
a = 8'd227; b = 8'd14;  #10 
a = 8'd227; b = 8'd15;  #10 
a = 8'd227; b = 8'd16;  #10 
a = 8'd227; b = 8'd17;  #10 
a = 8'd227; b = 8'd18;  #10 
a = 8'd227; b = 8'd19;  #10 
a = 8'd227; b = 8'd20;  #10 
a = 8'd227; b = 8'd21;  #10 
a = 8'd227; b = 8'd22;  #10 
a = 8'd227; b = 8'd23;  #10 
a = 8'd227; b = 8'd24;  #10 
a = 8'd227; b = 8'd25;  #10 
a = 8'd227; b = 8'd26;  #10 
a = 8'd227; b = 8'd27;  #10 
a = 8'd227; b = 8'd28;  #10 
a = 8'd227; b = 8'd29;  #10 
a = 8'd227; b = 8'd30;  #10 
a = 8'd227; b = 8'd31;  #10 
a = 8'd227; b = 8'd32;  #10 
a = 8'd227; b = 8'd33;  #10 
a = 8'd227; b = 8'd34;  #10 
a = 8'd227; b = 8'd35;  #10 
a = 8'd227; b = 8'd36;  #10 
a = 8'd227; b = 8'd37;  #10 
a = 8'd227; b = 8'd38;  #10 
a = 8'd227; b = 8'd39;  #10 
a = 8'd227; b = 8'd40;  #10 
a = 8'd227; b = 8'd41;  #10 
a = 8'd227; b = 8'd42;  #10 
a = 8'd227; b = 8'd43;  #10 
a = 8'd227; b = 8'd44;  #10 
a = 8'd227; b = 8'd45;  #10 
a = 8'd227; b = 8'd46;  #10 
a = 8'd227; b = 8'd47;  #10 
a = 8'd227; b = 8'd48;  #10 
a = 8'd227; b = 8'd49;  #10 
a = 8'd227; b = 8'd50;  #10 
a = 8'd227; b = 8'd51;  #10 
a = 8'd227; b = 8'd52;  #10 
a = 8'd227; b = 8'd53;  #10 
a = 8'd227; b = 8'd54;  #10 
a = 8'd227; b = 8'd55;  #10 
a = 8'd227; b = 8'd56;  #10 
a = 8'd227; b = 8'd57;  #10 
a = 8'd227; b = 8'd58;  #10 
a = 8'd227; b = 8'd59;  #10 
a = 8'd227; b = 8'd60;  #10 
a = 8'd227; b = 8'd61;  #10 
a = 8'd227; b = 8'd62;  #10 
a = 8'd227; b = 8'd63;  #10 
a = 8'd227; b = 8'd64;  #10 
a = 8'd227; b = 8'd65;  #10 
a = 8'd227; b = 8'd66;  #10 
a = 8'd227; b = 8'd67;  #10 
a = 8'd227; b = 8'd68;  #10 
a = 8'd227; b = 8'd69;  #10 
a = 8'd227; b = 8'd70;  #10 
a = 8'd227; b = 8'd71;  #10 
a = 8'd227; b = 8'd72;  #10 
a = 8'd227; b = 8'd73;  #10 
a = 8'd227; b = 8'd74;  #10 
a = 8'd227; b = 8'd75;  #10 
a = 8'd227; b = 8'd76;  #10 
a = 8'd227; b = 8'd77;  #10 
a = 8'd227; b = 8'd78;  #10 
a = 8'd227; b = 8'd79;  #10 
a = 8'd227; b = 8'd80;  #10 
a = 8'd227; b = 8'd81;  #10 
a = 8'd227; b = 8'd82;  #10 
a = 8'd227; b = 8'd83;  #10 
a = 8'd227; b = 8'd84;  #10 
a = 8'd227; b = 8'd85;  #10 
a = 8'd227; b = 8'd86;  #10 
a = 8'd227; b = 8'd87;  #10 
a = 8'd227; b = 8'd88;  #10 
a = 8'd227; b = 8'd89;  #10 
a = 8'd227; b = 8'd90;  #10 
a = 8'd227; b = 8'd91;  #10 
a = 8'd227; b = 8'd92;  #10 
a = 8'd227; b = 8'd93;  #10 
a = 8'd227; b = 8'd94;  #10 
a = 8'd227; b = 8'd95;  #10 
a = 8'd227; b = 8'd96;  #10 
a = 8'd227; b = 8'd97;  #10 
a = 8'd227; b = 8'd98;  #10 
a = 8'd227; b = 8'd99;  #10 
a = 8'd227; b = 8'd100;  #10 
a = 8'd227; b = 8'd101;  #10 
a = 8'd227; b = 8'd102;  #10 
a = 8'd227; b = 8'd103;  #10 
a = 8'd227; b = 8'd104;  #10 
a = 8'd227; b = 8'd105;  #10 
a = 8'd227; b = 8'd106;  #10 
a = 8'd227; b = 8'd107;  #10 
a = 8'd227; b = 8'd108;  #10 
a = 8'd227; b = 8'd109;  #10 
a = 8'd227; b = 8'd110;  #10 
a = 8'd227; b = 8'd111;  #10 
a = 8'd227; b = 8'd112;  #10 
a = 8'd227; b = 8'd113;  #10 
a = 8'd227; b = 8'd114;  #10 
a = 8'd227; b = 8'd115;  #10 
a = 8'd227; b = 8'd116;  #10 
a = 8'd227; b = 8'd117;  #10 
a = 8'd227; b = 8'd118;  #10 
a = 8'd227; b = 8'd119;  #10 
a = 8'd227; b = 8'd120;  #10 
a = 8'd227; b = 8'd121;  #10 
a = 8'd227; b = 8'd122;  #10 
a = 8'd227; b = 8'd123;  #10 
a = 8'd227; b = 8'd124;  #10 
a = 8'd227; b = 8'd125;  #10 
a = 8'd227; b = 8'd126;  #10 
a = 8'd227; b = 8'd127;  #10 
a = 8'd227; b = 8'd128;  #10 
a = 8'd227; b = 8'd129;  #10 
a = 8'd227; b = 8'd130;  #10 
a = 8'd227; b = 8'd131;  #10 
a = 8'd227; b = 8'd132;  #10 
a = 8'd227; b = 8'd133;  #10 
a = 8'd227; b = 8'd134;  #10 
a = 8'd227; b = 8'd135;  #10 
a = 8'd227; b = 8'd136;  #10 
a = 8'd227; b = 8'd137;  #10 
a = 8'd227; b = 8'd138;  #10 
a = 8'd227; b = 8'd139;  #10 
a = 8'd227; b = 8'd140;  #10 
a = 8'd227; b = 8'd141;  #10 
a = 8'd227; b = 8'd142;  #10 
a = 8'd227; b = 8'd143;  #10 
a = 8'd227; b = 8'd144;  #10 
a = 8'd227; b = 8'd145;  #10 
a = 8'd227; b = 8'd146;  #10 
a = 8'd227; b = 8'd147;  #10 
a = 8'd227; b = 8'd148;  #10 
a = 8'd227; b = 8'd149;  #10 
a = 8'd227; b = 8'd150;  #10 
a = 8'd227; b = 8'd151;  #10 
a = 8'd227; b = 8'd152;  #10 
a = 8'd227; b = 8'd153;  #10 
a = 8'd227; b = 8'd154;  #10 
a = 8'd227; b = 8'd155;  #10 
a = 8'd227; b = 8'd156;  #10 
a = 8'd227; b = 8'd157;  #10 
a = 8'd227; b = 8'd158;  #10 
a = 8'd227; b = 8'd159;  #10 
a = 8'd227; b = 8'd160;  #10 
a = 8'd227; b = 8'd161;  #10 
a = 8'd227; b = 8'd162;  #10 
a = 8'd227; b = 8'd163;  #10 
a = 8'd227; b = 8'd164;  #10 
a = 8'd227; b = 8'd165;  #10 
a = 8'd227; b = 8'd166;  #10 
a = 8'd227; b = 8'd167;  #10 
a = 8'd227; b = 8'd168;  #10 
a = 8'd227; b = 8'd169;  #10 
a = 8'd227; b = 8'd170;  #10 
a = 8'd227; b = 8'd171;  #10 
a = 8'd227; b = 8'd172;  #10 
a = 8'd227; b = 8'd173;  #10 
a = 8'd227; b = 8'd174;  #10 
a = 8'd227; b = 8'd175;  #10 
a = 8'd227; b = 8'd176;  #10 
a = 8'd227; b = 8'd177;  #10 
a = 8'd227; b = 8'd178;  #10 
a = 8'd227; b = 8'd179;  #10 
a = 8'd227; b = 8'd180;  #10 
a = 8'd227; b = 8'd181;  #10 
a = 8'd227; b = 8'd182;  #10 
a = 8'd227; b = 8'd183;  #10 
a = 8'd227; b = 8'd184;  #10 
a = 8'd227; b = 8'd185;  #10 
a = 8'd227; b = 8'd186;  #10 
a = 8'd227; b = 8'd187;  #10 
a = 8'd227; b = 8'd188;  #10 
a = 8'd227; b = 8'd189;  #10 
a = 8'd227; b = 8'd190;  #10 
a = 8'd227; b = 8'd191;  #10 
a = 8'd227; b = 8'd192;  #10 
a = 8'd227; b = 8'd193;  #10 
a = 8'd227; b = 8'd194;  #10 
a = 8'd227; b = 8'd195;  #10 
a = 8'd227; b = 8'd196;  #10 
a = 8'd227; b = 8'd197;  #10 
a = 8'd227; b = 8'd198;  #10 
a = 8'd227; b = 8'd199;  #10 
a = 8'd227; b = 8'd200;  #10 
a = 8'd227; b = 8'd201;  #10 
a = 8'd227; b = 8'd202;  #10 
a = 8'd227; b = 8'd203;  #10 
a = 8'd227; b = 8'd204;  #10 
a = 8'd227; b = 8'd205;  #10 
a = 8'd227; b = 8'd206;  #10 
a = 8'd227; b = 8'd207;  #10 
a = 8'd227; b = 8'd208;  #10 
a = 8'd227; b = 8'd209;  #10 
a = 8'd227; b = 8'd210;  #10 
a = 8'd227; b = 8'd211;  #10 
a = 8'd227; b = 8'd212;  #10 
a = 8'd227; b = 8'd213;  #10 
a = 8'd227; b = 8'd214;  #10 
a = 8'd227; b = 8'd215;  #10 
a = 8'd227; b = 8'd216;  #10 
a = 8'd227; b = 8'd217;  #10 
a = 8'd227; b = 8'd218;  #10 
a = 8'd227; b = 8'd219;  #10 
a = 8'd227; b = 8'd220;  #10 
a = 8'd227; b = 8'd221;  #10 
a = 8'd227; b = 8'd222;  #10 
a = 8'd227; b = 8'd223;  #10 
a = 8'd227; b = 8'd224;  #10 
a = 8'd227; b = 8'd225;  #10 
a = 8'd227; b = 8'd226;  #10 
a = 8'd227; b = 8'd227;  #10 
a = 8'd227; b = 8'd228;  #10 
a = 8'd227; b = 8'd229;  #10 
a = 8'd227; b = 8'd230;  #10 
a = 8'd227; b = 8'd231;  #10 
a = 8'd227; b = 8'd232;  #10 
a = 8'd227; b = 8'd233;  #10 
a = 8'd227; b = 8'd234;  #10 
a = 8'd227; b = 8'd235;  #10 
a = 8'd227; b = 8'd236;  #10 
a = 8'd227; b = 8'd237;  #10 
a = 8'd227; b = 8'd238;  #10 
a = 8'd227; b = 8'd239;  #10 
a = 8'd227; b = 8'd240;  #10 
a = 8'd227; b = 8'd241;  #10 
a = 8'd227; b = 8'd242;  #10 
a = 8'd227; b = 8'd243;  #10 
a = 8'd227; b = 8'd244;  #10 
a = 8'd227; b = 8'd245;  #10 
a = 8'd227; b = 8'd246;  #10 
a = 8'd227; b = 8'd247;  #10 
a = 8'd227; b = 8'd248;  #10 
a = 8'd227; b = 8'd249;  #10 
a = 8'd227; b = 8'd250;  #10 
a = 8'd227; b = 8'd251;  #10 
a = 8'd227; b = 8'd252;  #10 
a = 8'd227; b = 8'd253;  #10 
a = 8'd227; b = 8'd254;  #10 
a = 8'd227; b = 8'd255;  #10 
a = 8'd228; b = 8'd0;  #10 
a = 8'd228; b = 8'd1;  #10 
a = 8'd228; b = 8'd2;  #10 
a = 8'd228; b = 8'd3;  #10 
a = 8'd228; b = 8'd4;  #10 
a = 8'd228; b = 8'd5;  #10 
a = 8'd228; b = 8'd6;  #10 
a = 8'd228; b = 8'd7;  #10 
a = 8'd228; b = 8'd8;  #10 
a = 8'd228; b = 8'd9;  #10 
a = 8'd228; b = 8'd10;  #10 
a = 8'd228; b = 8'd11;  #10 
a = 8'd228; b = 8'd12;  #10 
a = 8'd228; b = 8'd13;  #10 
a = 8'd228; b = 8'd14;  #10 
a = 8'd228; b = 8'd15;  #10 
a = 8'd228; b = 8'd16;  #10 
a = 8'd228; b = 8'd17;  #10 
a = 8'd228; b = 8'd18;  #10 
a = 8'd228; b = 8'd19;  #10 
a = 8'd228; b = 8'd20;  #10 
a = 8'd228; b = 8'd21;  #10 
a = 8'd228; b = 8'd22;  #10 
a = 8'd228; b = 8'd23;  #10 
a = 8'd228; b = 8'd24;  #10 
a = 8'd228; b = 8'd25;  #10 
a = 8'd228; b = 8'd26;  #10 
a = 8'd228; b = 8'd27;  #10 
a = 8'd228; b = 8'd28;  #10 
a = 8'd228; b = 8'd29;  #10 
a = 8'd228; b = 8'd30;  #10 
a = 8'd228; b = 8'd31;  #10 
a = 8'd228; b = 8'd32;  #10 
a = 8'd228; b = 8'd33;  #10 
a = 8'd228; b = 8'd34;  #10 
a = 8'd228; b = 8'd35;  #10 
a = 8'd228; b = 8'd36;  #10 
a = 8'd228; b = 8'd37;  #10 
a = 8'd228; b = 8'd38;  #10 
a = 8'd228; b = 8'd39;  #10 
a = 8'd228; b = 8'd40;  #10 
a = 8'd228; b = 8'd41;  #10 
a = 8'd228; b = 8'd42;  #10 
a = 8'd228; b = 8'd43;  #10 
a = 8'd228; b = 8'd44;  #10 
a = 8'd228; b = 8'd45;  #10 
a = 8'd228; b = 8'd46;  #10 
a = 8'd228; b = 8'd47;  #10 
a = 8'd228; b = 8'd48;  #10 
a = 8'd228; b = 8'd49;  #10 
a = 8'd228; b = 8'd50;  #10 
a = 8'd228; b = 8'd51;  #10 
a = 8'd228; b = 8'd52;  #10 
a = 8'd228; b = 8'd53;  #10 
a = 8'd228; b = 8'd54;  #10 
a = 8'd228; b = 8'd55;  #10 
a = 8'd228; b = 8'd56;  #10 
a = 8'd228; b = 8'd57;  #10 
a = 8'd228; b = 8'd58;  #10 
a = 8'd228; b = 8'd59;  #10 
a = 8'd228; b = 8'd60;  #10 
a = 8'd228; b = 8'd61;  #10 
a = 8'd228; b = 8'd62;  #10 
a = 8'd228; b = 8'd63;  #10 
a = 8'd228; b = 8'd64;  #10 
a = 8'd228; b = 8'd65;  #10 
a = 8'd228; b = 8'd66;  #10 
a = 8'd228; b = 8'd67;  #10 
a = 8'd228; b = 8'd68;  #10 
a = 8'd228; b = 8'd69;  #10 
a = 8'd228; b = 8'd70;  #10 
a = 8'd228; b = 8'd71;  #10 
a = 8'd228; b = 8'd72;  #10 
a = 8'd228; b = 8'd73;  #10 
a = 8'd228; b = 8'd74;  #10 
a = 8'd228; b = 8'd75;  #10 
a = 8'd228; b = 8'd76;  #10 
a = 8'd228; b = 8'd77;  #10 
a = 8'd228; b = 8'd78;  #10 
a = 8'd228; b = 8'd79;  #10 
a = 8'd228; b = 8'd80;  #10 
a = 8'd228; b = 8'd81;  #10 
a = 8'd228; b = 8'd82;  #10 
a = 8'd228; b = 8'd83;  #10 
a = 8'd228; b = 8'd84;  #10 
a = 8'd228; b = 8'd85;  #10 
a = 8'd228; b = 8'd86;  #10 
a = 8'd228; b = 8'd87;  #10 
a = 8'd228; b = 8'd88;  #10 
a = 8'd228; b = 8'd89;  #10 
a = 8'd228; b = 8'd90;  #10 
a = 8'd228; b = 8'd91;  #10 
a = 8'd228; b = 8'd92;  #10 
a = 8'd228; b = 8'd93;  #10 
a = 8'd228; b = 8'd94;  #10 
a = 8'd228; b = 8'd95;  #10 
a = 8'd228; b = 8'd96;  #10 
a = 8'd228; b = 8'd97;  #10 
a = 8'd228; b = 8'd98;  #10 
a = 8'd228; b = 8'd99;  #10 
a = 8'd228; b = 8'd100;  #10 
a = 8'd228; b = 8'd101;  #10 
a = 8'd228; b = 8'd102;  #10 
a = 8'd228; b = 8'd103;  #10 
a = 8'd228; b = 8'd104;  #10 
a = 8'd228; b = 8'd105;  #10 
a = 8'd228; b = 8'd106;  #10 
a = 8'd228; b = 8'd107;  #10 
a = 8'd228; b = 8'd108;  #10 
a = 8'd228; b = 8'd109;  #10 
a = 8'd228; b = 8'd110;  #10 
a = 8'd228; b = 8'd111;  #10 
a = 8'd228; b = 8'd112;  #10 
a = 8'd228; b = 8'd113;  #10 
a = 8'd228; b = 8'd114;  #10 
a = 8'd228; b = 8'd115;  #10 
a = 8'd228; b = 8'd116;  #10 
a = 8'd228; b = 8'd117;  #10 
a = 8'd228; b = 8'd118;  #10 
a = 8'd228; b = 8'd119;  #10 
a = 8'd228; b = 8'd120;  #10 
a = 8'd228; b = 8'd121;  #10 
a = 8'd228; b = 8'd122;  #10 
a = 8'd228; b = 8'd123;  #10 
a = 8'd228; b = 8'd124;  #10 
a = 8'd228; b = 8'd125;  #10 
a = 8'd228; b = 8'd126;  #10 
a = 8'd228; b = 8'd127;  #10 
a = 8'd228; b = 8'd128;  #10 
a = 8'd228; b = 8'd129;  #10 
a = 8'd228; b = 8'd130;  #10 
a = 8'd228; b = 8'd131;  #10 
a = 8'd228; b = 8'd132;  #10 
a = 8'd228; b = 8'd133;  #10 
a = 8'd228; b = 8'd134;  #10 
a = 8'd228; b = 8'd135;  #10 
a = 8'd228; b = 8'd136;  #10 
a = 8'd228; b = 8'd137;  #10 
a = 8'd228; b = 8'd138;  #10 
a = 8'd228; b = 8'd139;  #10 
a = 8'd228; b = 8'd140;  #10 
a = 8'd228; b = 8'd141;  #10 
a = 8'd228; b = 8'd142;  #10 
a = 8'd228; b = 8'd143;  #10 
a = 8'd228; b = 8'd144;  #10 
a = 8'd228; b = 8'd145;  #10 
a = 8'd228; b = 8'd146;  #10 
a = 8'd228; b = 8'd147;  #10 
a = 8'd228; b = 8'd148;  #10 
a = 8'd228; b = 8'd149;  #10 
a = 8'd228; b = 8'd150;  #10 
a = 8'd228; b = 8'd151;  #10 
a = 8'd228; b = 8'd152;  #10 
a = 8'd228; b = 8'd153;  #10 
a = 8'd228; b = 8'd154;  #10 
a = 8'd228; b = 8'd155;  #10 
a = 8'd228; b = 8'd156;  #10 
a = 8'd228; b = 8'd157;  #10 
a = 8'd228; b = 8'd158;  #10 
a = 8'd228; b = 8'd159;  #10 
a = 8'd228; b = 8'd160;  #10 
a = 8'd228; b = 8'd161;  #10 
a = 8'd228; b = 8'd162;  #10 
a = 8'd228; b = 8'd163;  #10 
a = 8'd228; b = 8'd164;  #10 
a = 8'd228; b = 8'd165;  #10 
a = 8'd228; b = 8'd166;  #10 
a = 8'd228; b = 8'd167;  #10 
a = 8'd228; b = 8'd168;  #10 
a = 8'd228; b = 8'd169;  #10 
a = 8'd228; b = 8'd170;  #10 
a = 8'd228; b = 8'd171;  #10 
a = 8'd228; b = 8'd172;  #10 
a = 8'd228; b = 8'd173;  #10 
a = 8'd228; b = 8'd174;  #10 
a = 8'd228; b = 8'd175;  #10 
a = 8'd228; b = 8'd176;  #10 
a = 8'd228; b = 8'd177;  #10 
a = 8'd228; b = 8'd178;  #10 
a = 8'd228; b = 8'd179;  #10 
a = 8'd228; b = 8'd180;  #10 
a = 8'd228; b = 8'd181;  #10 
a = 8'd228; b = 8'd182;  #10 
a = 8'd228; b = 8'd183;  #10 
a = 8'd228; b = 8'd184;  #10 
a = 8'd228; b = 8'd185;  #10 
a = 8'd228; b = 8'd186;  #10 
a = 8'd228; b = 8'd187;  #10 
a = 8'd228; b = 8'd188;  #10 
a = 8'd228; b = 8'd189;  #10 
a = 8'd228; b = 8'd190;  #10 
a = 8'd228; b = 8'd191;  #10 
a = 8'd228; b = 8'd192;  #10 
a = 8'd228; b = 8'd193;  #10 
a = 8'd228; b = 8'd194;  #10 
a = 8'd228; b = 8'd195;  #10 
a = 8'd228; b = 8'd196;  #10 
a = 8'd228; b = 8'd197;  #10 
a = 8'd228; b = 8'd198;  #10 
a = 8'd228; b = 8'd199;  #10 
a = 8'd228; b = 8'd200;  #10 
a = 8'd228; b = 8'd201;  #10 
a = 8'd228; b = 8'd202;  #10 
a = 8'd228; b = 8'd203;  #10 
a = 8'd228; b = 8'd204;  #10 
a = 8'd228; b = 8'd205;  #10 
a = 8'd228; b = 8'd206;  #10 
a = 8'd228; b = 8'd207;  #10 
a = 8'd228; b = 8'd208;  #10 
a = 8'd228; b = 8'd209;  #10 
a = 8'd228; b = 8'd210;  #10 
a = 8'd228; b = 8'd211;  #10 
a = 8'd228; b = 8'd212;  #10 
a = 8'd228; b = 8'd213;  #10 
a = 8'd228; b = 8'd214;  #10 
a = 8'd228; b = 8'd215;  #10 
a = 8'd228; b = 8'd216;  #10 
a = 8'd228; b = 8'd217;  #10 
a = 8'd228; b = 8'd218;  #10 
a = 8'd228; b = 8'd219;  #10 
a = 8'd228; b = 8'd220;  #10 
a = 8'd228; b = 8'd221;  #10 
a = 8'd228; b = 8'd222;  #10 
a = 8'd228; b = 8'd223;  #10 
a = 8'd228; b = 8'd224;  #10 
a = 8'd228; b = 8'd225;  #10 
a = 8'd228; b = 8'd226;  #10 
a = 8'd228; b = 8'd227;  #10 
a = 8'd228; b = 8'd228;  #10 
a = 8'd228; b = 8'd229;  #10 
a = 8'd228; b = 8'd230;  #10 
a = 8'd228; b = 8'd231;  #10 
a = 8'd228; b = 8'd232;  #10 
a = 8'd228; b = 8'd233;  #10 
a = 8'd228; b = 8'd234;  #10 
a = 8'd228; b = 8'd235;  #10 
a = 8'd228; b = 8'd236;  #10 
a = 8'd228; b = 8'd237;  #10 
a = 8'd228; b = 8'd238;  #10 
a = 8'd228; b = 8'd239;  #10 
a = 8'd228; b = 8'd240;  #10 
a = 8'd228; b = 8'd241;  #10 
a = 8'd228; b = 8'd242;  #10 
a = 8'd228; b = 8'd243;  #10 
a = 8'd228; b = 8'd244;  #10 
a = 8'd228; b = 8'd245;  #10 
a = 8'd228; b = 8'd246;  #10 
a = 8'd228; b = 8'd247;  #10 
a = 8'd228; b = 8'd248;  #10 
a = 8'd228; b = 8'd249;  #10 
a = 8'd228; b = 8'd250;  #10 
a = 8'd228; b = 8'd251;  #10 
a = 8'd228; b = 8'd252;  #10 
a = 8'd228; b = 8'd253;  #10 
a = 8'd228; b = 8'd254;  #10 
a = 8'd228; b = 8'd255;  #10 
a = 8'd229; b = 8'd0;  #10 
a = 8'd229; b = 8'd1;  #10 
a = 8'd229; b = 8'd2;  #10 
a = 8'd229; b = 8'd3;  #10 
a = 8'd229; b = 8'd4;  #10 
a = 8'd229; b = 8'd5;  #10 
a = 8'd229; b = 8'd6;  #10 
a = 8'd229; b = 8'd7;  #10 
a = 8'd229; b = 8'd8;  #10 
a = 8'd229; b = 8'd9;  #10 
a = 8'd229; b = 8'd10;  #10 
a = 8'd229; b = 8'd11;  #10 
a = 8'd229; b = 8'd12;  #10 
a = 8'd229; b = 8'd13;  #10 
a = 8'd229; b = 8'd14;  #10 
a = 8'd229; b = 8'd15;  #10 
a = 8'd229; b = 8'd16;  #10 
a = 8'd229; b = 8'd17;  #10 
a = 8'd229; b = 8'd18;  #10 
a = 8'd229; b = 8'd19;  #10 
a = 8'd229; b = 8'd20;  #10 
a = 8'd229; b = 8'd21;  #10 
a = 8'd229; b = 8'd22;  #10 
a = 8'd229; b = 8'd23;  #10 
a = 8'd229; b = 8'd24;  #10 
a = 8'd229; b = 8'd25;  #10 
a = 8'd229; b = 8'd26;  #10 
a = 8'd229; b = 8'd27;  #10 
a = 8'd229; b = 8'd28;  #10 
a = 8'd229; b = 8'd29;  #10 
a = 8'd229; b = 8'd30;  #10 
a = 8'd229; b = 8'd31;  #10 
a = 8'd229; b = 8'd32;  #10 
a = 8'd229; b = 8'd33;  #10 
a = 8'd229; b = 8'd34;  #10 
a = 8'd229; b = 8'd35;  #10 
a = 8'd229; b = 8'd36;  #10 
a = 8'd229; b = 8'd37;  #10 
a = 8'd229; b = 8'd38;  #10 
a = 8'd229; b = 8'd39;  #10 
a = 8'd229; b = 8'd40;  #10 
a = 8'd229; b = 8'd41;  #10 
a = 8'd229; b = 8'd42;  #10 
a = 8'd229; b = 8'd43;  #10 
a = 8'd229; b = 8'd44;  #10 
a = 8'd229; b = 8'd45;  #10 
a = 8'd229; b = 8'd46;  #10 
a = 8'd229; b = 8'd47;  #10 
a = 8'd229; b = 8'd48;  #10 
a = 8'd229; b = 8'd49;  #10 
a = 8'd229; b = 8'd50;  #10 
a = 8'd229; b = 8'd51;  #10 
a = 8'd229; b = 8'd52;  #10 
a = 8'd229; b = 8'd53;  #10 
a = 8'd229; b = 8'd54;  #10 
a = 8'd229; b = 8'd55;  #10 
a = 8'd229; b = 8'd56;  #10 
a = 8'd229; b = 8'd57;  #10 
a = 8'd229; b = 8'd58;  #10 
a = 8'd229; b = 8'd59;  #10 
a = 8'd229; b = 8'd60;  #10 
a = 8'd229; b = 8'd61;  #10 
a = 8'd229; b = 8'd62;  #10 
a = 8'd229; b = 8'd63;  #10 
a = 8'd229; b = 8'd64;  #10 
a = 8'd229; b = 8'd65;  #10 
a = 8'd229; b = 8'd66;  #10 
a = 8'd229; b = 8'd67;  #10 
a = 8'd229; b = 8'd68;  #10 
a = 8'd229; b = 8'd69;  #10 
a = 8'd229; b = 8'd70;  #10 
a = 8'd229; b = 8'd71;  #10 
a = 8'd229; b = 8'd72;  #10 
a = 8'd229; b = 8'd73;  #10 
a = 8'd229; b = 8'd74;  #10 
a = 8'd229; b = 8'd75;  #10 
a = 8'd229; b = 8'd76;  #10 
a = 8'd229; b = 8'd77;  #10 
a = 8'd229; b = 8'd78;  #10 
a = 8'd229; b = 8'd79;  #10 
a = 8'd229; b = 8'd80;  #10 
a = 8'd229; b = 8'd81;  #10 
a = 8'd229; b = 8'd82;  #10 
a = 8'd229; b = 8'd83;  #10 
a = 8'd229; b = 8'd84;  #10 
a = 8'd229; b = 8'd85;  #10 
a = 8'd229; b = 8'd86;  #10 
a = 8'd229; b = 8'd87;  #10 
a = 8'd229; b = 8'd88;  #10 
a = 8'd229; b = 8'd89;  #10 
a = 8'd229; b = 8'd90;  #10 
a = 8'd229; b = 8'd91;  #10 
a = 8'd229; b = 8'd92;  #10 
a = 8'd229; b = 8'd93;  #10 
a = 8'd229; b = 8'd94;  #10 
a = 8'd229; b = 8'd95;  #10 
a = 8'd229; b = 8'd96;  #10 
a = 8'd229; b = 8'd97;  #10 
a = 8'd229; b = 8'd98;  #10 
a = 8'd229; b = 8'd99;  #10 
a = 8'd229; b = 8'd100;  #10 
a = 8'd229; b = 8'd101;  #10 
a = 8'd229; b = 8'd102;  #10 
a = 8'd229; b = 8'd103;  #10 
a = 8'd229; b = 8'd104;  #10 
a = 8'd229; b = 8'd105;  #10 
a = 8'd229; b = 8'd106;  #10 
a = 8'd229; b = 8'd107;  #10 
a = 8'd229; b = 8'd108;  #10 
a = 8'd229; b = 8'd109;  #10 
a = 8'd229; b = 8'd110;  #10 
a = 8'd229; b = 8'd111;  #10 
a = 8'd229; b = 8'd112;  #10 
a = 8'd229; b = 8'd113;  #10 
a = 8'd229; b = 8'd114;  #10 
a = 8'd229; b = 8'd115;  #10 
a = 8'd229; b = 8'd116;  #10 
a = 8'd229; b = 8'd117;  #10 
a = 8'd229; b = 8'd118;  #10 
a = 8'd229; b = 8'd119;  #10 
a = 8'd229; b = 8'd120;  #10 
a = 8'd229; b = 8'd121;  #10 
a = 8'd229; b = 8'd122;  #10 
a = 8'd229; b = 8'd123;  #10 
a = 8'd229; b = 8'd124;  #10 
a = 8'd229; b = 8'd125;  #10 
a = 8'd229; b = 8'd126;  #10 
a = 8'd229; b = 8'd127;  #10 
a = 8'd229; b = 8'd128;  #10 
a = 8'd229; b = 8'd129;  #10 
a = 8'd229; b = 8'd130;  #10 
a = 8'd229; b = 8'd131;  #10 
a = 8'd229; b = 8'd132;  #10 
a = 8'd229; b = 8'd133;  #10 
a = 8'd229; b = 8'd134;  #10 
a = 8'd229; b = 8'd135;  #10 
a = 8'd229; b = 8'd136;  #10 
a = 8'd229; b = 8'd137;  #10 
a = 8'd229; b = 8'd138;  #10 
a = 8'd229; b = 8'd139;  #10 
a = 8'd229; b = 8'd140;  #10 
a = 8'd229; b = 8'd141;  #10 
a = 8'd229; b = 8'd142;  #10 
a = 8'd229; b = 8'd143;  #10 
a = 8'd229; b = 8'd144;  #10 
a = 8'd229; b = 8'd145;  #10 
a = 8'd229; b = 8'd146;  #10 
a = 8'd229; b = 8'd147;  #10 
a = 8'd229; b = 8'd148;  #10 
a = 8'd229; b = 8'd149;  #10 
a = 8'd229; b = 8'd150;  #10 
a = 8'd229; b = 8'd151;  #10 
a = 8'd229; b = 8'd152;  #10 
a = 8'd229; b = 8'd153;  #10 
a = 8'd229; b = 8'd154;  #10 
a = 8'd229; b = 8'd155;  #10 
a = 8'd229; b = 8'd156;  #10 
a = 8'd229; b = 8'd157;  #10 
a = 8'd229; b = 8'd158;  #10 
a = 8'd229; b = 8'd159;  #10 
a = 8'd229; b = 8'd160;  #10 
a = 8'd229; b = 8'd161;  #10 
a = 8'd229; b = 8'd162;  #10 
a = 8'd229; b = 8'd163;  #10 
a = 8'd229; b = 8'd164;  #10 
a = 8'd229; b = 8'd165;  #10 
a = 8'd229; b = 8'd166;  #10 
a = 8'd229; b = 8'd167;  #10 
a = 8'd229; b = 8'd168;  #10 
a = 8'd229; b = 8'd169;  #10 
a = 8'd229; b = 8'd170;  #10 
a = 8'd229; b = 8'd171;  #10 
a = 8'd229; b = 8'd172;  #10 
a = 8'd229; b = 8'd173;  #10 
a = 8'd229; b = 8'd174;  #10 
a = 8'd229; b = 8'd175;  #10 
a = 8'd229; b = 8'd176;  #10 
a = 8'd229; b = 8'd177;  #10 
a = 8'd229; b = 8'd178;  #10 
a = 8'd229; b = 8'd179;  #10 
a = 8'd229; b = 8'd180;  #10 
a = 8'd229; b = 8'd181;  #10 
a = 8'd229; b = 8'd182;  #10 
a = 8'd229; b = 8'd183;  #10 
a = 8'd229; b = 8'd184;  #10 
a = 8'd229; b = 8'd185;  #10 
a = 8'd229; b = 8'd186;  #10 
a = 8'd229; b = 8'd187;  #10 
a = 8'd229; b = 8'd188;  #10 
a = 8'd229; b = 8'd189;  #10 
a = 8'd229; b = 8'd190;  #10 
a = 8'd229; b = 8'd191;  #10 
a = 8'd229; b = 8'd192;  #10 
a = 8'd229; b = 8'd193;  #10 
a = 8'd229; b = 8'd194;  #10 
a = 8'd229; b = 8'd195;  #10 
a = 8'd229; b = 8'd196;  #10 
a = 8'd229; b = 8'd197;  #10 
a = 8'd229; b = 8'd198;  #10 
a = 8'd229; b = 8'd199;  #10 
a = 8'd229; b = 8'd200;  #10 
a = 8'd229; b = 8'd201;  #10 
a = 8'd229; b = 8'd202;  #10 
a = 8'd229; b = 8'd203;  #10 
a = 8'd229; b = 8'd204;  #10 
a = 8'd229; b = 8'd205;  #10 
a = 8'd229; b = 8'd206;  #10 
a = 8'd229; b = 8'd207;  #10 
a = 8'd229; b = 8'd208;  #10 
a = 8'd229; b = 8'd209;  #10 
a = 8'd229; b = 8'd210;  #10 
a = 8'd229; b = 8'd211;  #10 
a = 8'd229; b = 8'd212;  #10 
a = 8'd229; b = 8'd213;  #10 
a = 8'd229; b = 8'd214;  #10 
a = 8'd229; b = 8'd215;  #10 
a = 8'd229; b = 8'd216;  #10 
a = 8'd229; b = 8'd217;  #10 
a = 8'd229; b = 8'd218;  #10 
a = 8'd229; b = 8'd219;  #10 
a = 8'd229; b = 8'd220;  #10 
a = 8'd229; b = 8'd221;  #10 
a = 8'd229; b = 8'd222;  #10 
a = 8'd229; b = 8'd223;  #10 
a = 8'd229; b = 8'd224;  #10 
a = 8'd229; b = 8'd225;  #10 
a = 8'd229; b = 8'd226;  #10 
a = 8'd229; b = 8'd227;  #10 
a = 8'd229; b = 8'd228;  #10 
a = 8'd229; b = 8'd229;  #10 
a = 8'd229; b = 8'd230;  #10 
a = 8'd229; b = 8'd231;  #10 
a = 8'd229; b = 8'd232;  #10 
a = 8'd229; b = 8'd233;  #10 
a = 8'd229; b = 8'd234;  #10 
a = 8'd229; b = 8'd235;  #10 
a = 8'd229; b = 8'd236;  #10 
a = 8'd229; b = 8'd237;  #10 
a = 8'd229; b = 8'd238;  #10 
a = 8'd229; b = 8'd239;  #10 
a = 8'd229; b = 8'd240;  #10 
a = 8'd229; b = 8'd241;  #10 
a = 8'd229; b = 8'd242;  #10 
a = 8'd229; b = 8'd243;  #10 
a = 8'd229; b = 8'd244;  #10 
a = 8'd229; b = 8'd245;  #10 
a = 8'd229; b = 8'd246;  #10 
a = 8'd229; b = 8'd247;  #10 
a = 8'd229; b = 8'd248;  #10 
a = 8'd229; b = 8'd249;  #10 
a = 8'd229; b = 8'd250;  #10 
a = 8'd229; b = 8'd251;  #10 
a = 8'd229; b = 8'd252;  #10 
a = 8'd229; b = 8'd253;  #10 
a = 8'd229; b = 8'd254;  #10 
a = 8'd229; b = 8'd255;  #10 
a = 8'd230; b = 8'd0;  #10 
a = 8'd230; b = 8'd1;  #10 
a = 8'd230; b = 8'd2;  #10 
a = 8'd230; b = 8'd3;  #10 
a = 8'd230; b = 8'd4;  #10 
a = 8'd230; b = 8'd5;  #10 
a = 8'd230; b = 8'd6;  #10 
a = 8'd230; b = 8'd7;  #10 
a = 8'd230; b = 8'd8;  #10 
a = 8'd230; b = 8'd9;  #10 
a = 8'd230; b = 8'd10;  #10 
a = 8'd230; b = 8'd11;  #10 
a = 8'd230; b = 8'd12;  #10 
a = 8'd230; b = 8'd13;  #10 
a = 8'd230; b = 8'd14;  #10 
a = 8'd230; b = 8'd15;  #10 
a = 8'd230; b = 8'd16;  #10 
a = 8'd230; b = 8'd17;  #10 
a = 8'd230; b = 8'd18;  #10 
a = 8'd230; b = 8'd19;  #10 
a = 8'd230; b = 8'd20;  #10 
a = 8'd230; b = 8'd21;  #10 
a = 8'd230; b = 8'd22;  #10 
a = 8'd230; b = 8'd23;  #10 
a = 8'd230; b = 8'd24;  #10 
a = 8'd230; b = 8'd25;  #10 
a = 8'd230; b = 8'd26;  #10 
a = 8'd230; b = 8'd27;  #10 
a = 8'd230; b = 8'd28;  #10 
a = 8'd230; b = 8'd29;  #10 
a = 8'd230; b = 8'd30;  #10 
a = 8'd230; b = 8'd31;  #10 
a = 8'd230; b = 8'd32;  #10 
a = 8'd230; b = 8'd33;  #10 
a = 8'd230; b = 8'd34;  #10 
a = 8'd230; b = 8'd35;  #10 
a = 8'd230; b = 8'd36;  #10 
a = 8'd230; b = 8'd37;  #10 
a = 8'd230; b = 8'd38;  #10 
a = 8'd230; b = 8'd39;  #10 
a = 8'd230; b = 8'd40;  #10 
a = 8'd230; b = 8'd41;  #10 
a = 8'd230; b = 8'd42;  #10 
a = 8'd230; b = 8'd43;  #10 
a = 8'd230; b = 8'd44;  #10 
a = 8'd230; b = 8'd45;  #10 
a = 8'd230; b = 8'd46;  #10 
a = 8'd230; b = 8'd47;  #10 
a = 8'd230; b = 8'd48;  #10 
a = 8'd230; b = 8'd49;  #10 
a = 8'd230; b = 8'd50;  #10 
a = 8'd230; b = 8'd51;  #10 
a = 8'd230; b = 8'd52;  #10 
a = 8'd230; b = 8'd53;  #10 
a = 8'd230; b = 8'd54;  #10 
a = 8'd230; b = 8'd55;  #10 
a = 8'd230; b = 8'd56;  #10 
a = 8'd230; b = 8'd57;  #10 
a = 8'd230; b = 8'd58;  #10 
a = 8'd230; b = 8'd59;  #10 
a = 8'd230; b = 8'd60;  #10 
a = 8'd230; b = 8'd61;  #10 
a = 8'd230; b = 8'd62;  #10 
a = 8'd230; b = 8'd63;  #10 
a = 8'd230; b = 8'd64;  #10 
a = 8'd230; b = 8'd65;  #10 
a = 8'd230; b = 8'd66;  #10 
a = 8'd230; b = 8'd67;  #10 
a = 8'd230; b = 8'd68;  #10 
a = 8'd230; b = 8'd69;  #10 
a = 8'd230; b = 8'd70;  #10 
a = 8'd230; b = 8'd71;  #10 
a = 8'd230; b = 8'd72;  #10 
a = 8'd230; b = 8'd73;  #10 
a = 8'd230; b = 8'd74;  #10 
a = 8'd230; b = 8'd75;  #10 
a = 8'd230; b = 8'd76;  #10 
a = 8'd230; b = 8'd77;  #10 
a = 8'd230; b = 8'd78;  #10 
a = 8'd230; b = 8'd79;  #10 
a = 8'd230; b = 8'd80;  #10 
a = 8'd230; b = 8'd81;  #10 
a = 8'd230; b = 8'd82;  #10 
a = 8'd230; b = 8'd83;  #10 
a = 8'd230; b = 8'd84;  #10 
a = 8'd230; b = 8'd85;  #10 
a = 8'd230; b = 8'd86;  #10 
a = 8'd230; b = 8'd87;  #10 
a = 8'd230; b = 8'd88;  #10 
a = 8'd230; b = 8'd89;  #10 
a = 8'd230; b = 8'd90;  #10 
a = 8'd230; b = 8'd91;  #10 
a = 8'd230; b = 8'd92;  #10 
a = 8'd230; b = 8'd93;  #10 
a = 8'd230; b = 8'd94;  #10 
a = 8'd230; b = 8'd95;  #10 
a = 8'd230; b = 8'd96;  #10 
a = 8'd230; b = 8'd97;  #10 
a = 8'd230; b = 8'd98;  #10 
a = 8'd230; b = 8'd99;  #10 
a = 8'd230; b = 8'd100;  #10 
a = 8'd230; b = 8'd101;  #10 
a = 8'd230; b = 8'd102;  #10 
a = 8'd230; b = 8'd103;  #10 
a = 8'd230; b = 8'd104;  #10 
a = 8'd230; b = 8'd105;  #10 
a = 8'd230; b = 8'd106;  #10 
a = 8'd230; b = 8'd107;  #10 
a = 8'd230; b = 8'd108;  #10 
a = 8'd230; b = 8'd109;  #10 
a = 8'd230; b = 8'd110;  #10 
a = 8'd230; b = 8'd111;  #10 
a = 8'd230; b = 8'd112;  #10 
a = 8'd230; b = 8'd113;  #10 
a = 8'd230; b = 8'd114;  #10 
a = 8'd230; b = 8'd115;  #10 
a = 8'd230; b = 8'd116;  #10 
a = 8'd230; b = 8'd117;  #10 
a = 8'd230; b = 8'd118;  #10 
a = 8'd230; b = 8'd119;  #10 
a = 8'd230; b = 8'd120;  #10 
a = 8'd230; b = 8'd121;  #10 
a = 8'd230; b = 8'd122;  #10 
a = 8'd230; b = 8'd123;  #10 
a = 8'd230; b = 8'd124;  #10 
a = 8'd230; b = 8'd125;  #10 
a = 8'd230; b = 8'd126;  #10 
a = 8'd230; b = 8'd127;  #10 
a = 8'd230; b = 8'd128;  #10 
a = 8'd230; b = 8'd129;  #10 
a = 8'd230; b = 8'd130;  #10 
a = 8'd230; b = 8'd131;  #10 
a = 8'd230; b = 8'd132;  #10 
a = 8'd230; b = 8'd133;  #10 
a = 8'd230; b = 8'd134;  #10 
a = 8'd230; b = 8'd135;  #10 
a = 8'd230; b = 8'd136;  #10 
a = 8'd230; b = 8'd137;  #10 
a = 8'd230; b = 8'd138;  #10 
a = 8'd230; b = 8'd139;  #10 
a = 8'd230; b = 8'd140;  #10 
a = 8'd230; b = 8'd141;  #10 
a = 8'd230; b = 8'd142;  #10 
a = 8'd230; b = 8'd143;  #10 
a = 8'd230; b = 8'd144;  #10 
a = 8'd230; b = 8'd145;  #10 
a = 8'd230; b = 8'd146;  #10 
a = 8'd230; b = 8'd147;  #10 
a = 8'd230; b = 8'd148;  #10 
a = 8'd230; b = 8'd149;  #10 
a = 8'd230; b = 8'd150;  #10 
a = 8'd230; b = 8'd151;  #10 
a = 8'd230; b = 8'd152;  #10 
a = 8'd230; b = 8'd153;  #10 
a = 8'd230; b = 8'd154;  #10 
a = 8'd230; b = 8'd155;  #10 
a = 8'd230; b = 8'd156;  #10 
a = 8'd230; b = 8'd157;  #10 
a = 8'd230; b = 8'd158;  #10 
a = 8'd230; b = 8'd159;  #10 
a = 8'd230; b = 8'd160;  #10 
a = 8'd230; b = 8'd161;  #10 
a = 8'd230; b = 8'd162;  #10 
a = 8'd230; b = 8'd163;  #10 
a = 8'd230; b = 8'd164;  #10 
a = 8'd230; b = 8'd165;  #10 
a = 8'd230; b = 8'd166;  #10 
a = 8'd230; b = 8'd167;  #10 
a = 8'd230; b = 8'd168;  #10 
a = 8'd230; b = 8'd169;  #10 
a = 8'd230; b = 8'd170;  #10 
a = 8'd230; b = 8'd171;  #10 
a = 8'd230; b = 8'd172;  #10 
a = 8'd230; b = 8'd173;  #10 
a = 8'd230; b = 8'd174;  #10 
a = 8'd230; b = 8'd175;  #10 
a = 8'd230; b = 8'd176;  #10 
a = 8'd230; b = 8'd177;  #10 
a = 8'd230; b = 8'd178;  #10 
a = 8'd230; b = 8'd179;  #10 
a = 8'd230; b = 8'd180;  #10 
a = 8'd230; b = 8'd181;  #10 
a = 8'd230; b = 8'd182;  #10 
a = 8'd230; b = 8'd183;  #10 
a = 8'd230; b = 8'd184;  #10 
a = 8'd230; b = 8'd185;  #10 
a = 8'd230; b = 8'd186;  #10 
a = 8'd230; b = 8'd187;  #10 
a = 8'd230; b = 8'd188;  #10 
a = 8'd230; b = 8'd189;  #10 
a = 8'd230; b = 8'd190;  #10 
a = 8'd230; b = 8'd191;  #10 
a = 8'd230; b = 8'd192;  #10 
a = 8'd230; b = 8'd193;  #10 
a = 8'd230; b = 8'd194;  #10 
a = 8'd230; b = 8'd195;  #10 
a = 8'd230; b = 8'd196;  #10 
a = 8'd230; b = 8'd197;  #10 
a = 8'd230; b = 8'd198;  #10 
a = 8'd230; b = 8'd199;  #10 
a = 8'd230; b = 8'd200;  #10 
a = 8'd230; b = 8'd201;  #10 
a = 8'd230; b = 8'd202;  #10 
a = 8'd230; b = 8'd203;  #10 
a = 8'd230; b = 8'd204;  #10 
a = 8'd230; b = 8'd205;  #10 
a = 8'd230; b = 8'd206;  #10 
a = 8'd230; b = 8'd207;  #10 
a = 8'd230; b = 8'd208;  #10 
a = 8'd230; b = 8'd209;  #10 
a = 8'd230; b = 8'd210;  #10 
a = 8'd230; b = 8'd211;  #10 
a = 8'd230; b = 8'd212;  #10 
a = 8'd230; b = 8'd213;  #10 
a = 8'd230; b = 8'd214;  #10 
a = 8'd230; b = 8'd215;  #10 
a = 8'd230; b = 8'd216;  #10 
a = 8'd230; b = 8'd217;  #10 
a = 8'd230; b = 8'd218;  #10 
a = 8'd230; b = 8'd219;  #10 
a = 8'd230; b = 8'd220;  #10 
a = 8'd230; b = 8'd221;  #10 
a = 8'd230; b = 8'd222;  #10 
a = 8'd230; b = 8'd223;  #10 
a = 8'd230; b = 8'd224;  #10 
a = 8'd230; b = 8'd225;  #10 
a = 8'd230; b = 8'd226;  #10 
a = 8'd230; b = 8'd227;  #10 
a = 8'd230; b = 8'd228;  #10 
a = 8'd230; b = 8'd229;  #10 
a = 8'd230; b = 8'd230;  #10 
a = 8'd230; b = 8'd231;  #10 
a = 8'd230; b = 8'd232;  #10 
a = 8'd230; b = 8'd233;  #10 
a = 8'd230; b = 8'd234;  #10 
a = 8'd230; b = 8'd235;  #10 
a = 8'd230; b = 8'd236;  #10 
a = 8'd230; b = 8'd237;  #10 
a = 8'd230; b = 8'd238;  #10 
a = 8'd230; b = 8'd239;  #10 
a = 8'd230; b = 8'd240;  #10 
a = 8'd230; b = 8'd241;  #10 
a = 8'd230; b = 8'd242;  #10 
a = 8'd230; b = 8'd243;  #10 
a = 8'd230; b = 8'd244;  #10 
a = 8'd230; b = 8'd245;  #10 
a = 8'd230; b = 8'd246;  #10 
a = 8'd230; b = 8'd247;  #10 
a = 8'd230; b = 8'd248;  #10 
a = 8'd230; b = 8'd249;  #10 
a = 8'd230; b = 8'd250;  #10 
a = 8'd230; b = 8'd251;  #10 
a = 8'd230; b = 8'd252;  #10 
a = 8'd230; b = 8'd253;  #10 
a = 8'd230; b = 8'd254;  #10 
a = 8'd230; b = 8'd255;  #10 
a = 8'd231; b = 8'd0;  #10 
a = 8'd231; b = 8'd1;  #10 
a = 8'd231; b = 8'd2;  #10 
a = 8'd231; b = 8'd3;  #10 
a = 8'd231; b = 8'd4;  #10 
a = 8'd231; b = 8'd5;  #10 
a = 8'd231; b = 8'd6;  #10 
a = 8'd231; b = 8'd7;  #10 
a = 8'd231; b = 8'd8;  #10 
a = 8'd231; b = 8'd9;  #10 
a = 8'd231; b = 8'd10;  #10 
a = 8'd231; b = 8'd11;  #10 
a = 8'd231; b = 8'd12;  #10 
a = 8'd231; b = 8'd13;  #10 
a = 8'd231; b = 8'd14;  #10 
a = 8'd231; b = 8'd15;  #10 
a = 8'd231; b = 8'd16;  #10 
a = 8'd231; b = 8'd17;  #10 
a = 8'd231; b = 8'd18;  #10 
a = 8'd231; b = 8'd19;  #10 
a = 8'd231; b = 8'd20;  #10 
a = 8'd231; b = 8'd21;  #10 
a = 8'd231; b = 8'd22;  #10 
a = 8'd231; b = 8'd23;  #10 
a = 8'd231; b = 8'd24;  #10 
a = 8'd231; b = 8'd25;  #10 
a = 8'd231; b = 8'd26;  #10 
a = 8'd231; b = 8'd27;  #10 
a = 8'd231; b = 8'd28;  #10 
a = 8'd231; b = 8'd29;  #10 
a = 8'd231; b = 8'd30;  #10 
a = 8'd231; b = 8'd31;  #10 
a = 8'd231; b = 8'd32;  #10 
a = 8'd231; b = 8'd33;  #10 
a = 8'd231; b = 8'd34;  #10 
a = 8'd231; b = 8'd35;  #10 
a = 8'd231; b = 8'd36;  #10 
a = 8'd231; b = 8'd37;  #10 
a = 8'd231; b = 8'd38;  #10 
a = 8'd231; b = 8'd39;  #10 
a = 8'd231; b = 8'd40;  #10 
a = 8'd231; b = 8'd41;  #10 
a = 8'd231; b = 8'd42;  #10 
a = 8'd231; b = 8'd43;  #10 
a = 8'd231; b = 8'd44;  #10 
a = 8'd231; b = 8'd45;  #10 
a = 8'd231; b = 8'd46;  #10 
a = 8'd231; b = 8'd47;  #10 
a = 8'd231; b = 8'd48;  #10 
a = 8'd231; b = 8'd49;  #10 
a = 8'd231; b = 8'd50;  #10 
a = 8'd231; b = 8'd51;  #10 
a = 8'd231; b = 8'd52;  #10 
a = 8'd231; b = 8'd53;  #10 
a = 8'd231; b = 8'd54;  #10 
a = 8'd231; b = 8'd55;  #10 
a = 8'd231; b = 8'd56;  #10 
a = 8'd231; b = 8'd57;  #10 
a = 8'd231; b = 8'd58;  #10 
a = 8'd231; b = 8'd59;  #10 
a = 8'd231; b = 8'd60;  #10 
a = 8'd231; b = 8'd61;  #10 
a = 8'd231; b = 8'd62;  #10 
a = 8'd231; b = 8'd63;  #10 
a = 8'd231; b = 8'd64;  #10 
a = 8'd231; b = 8'd65;  #10 
a = 8'd231; b = 8'd66;  #10 
a = 8'd231; b = 8'd67;  #10 
a = 8'd231; b = 8'd68;  #10 
a = 8'd231; b = 8'd69;  #10 
a = 8'd231; b = 8'd70;  #10 
a = 8'd231; b = 8'd71;  #10 
a = 8'd231; b = 8'd72;  #10 
a = 8'd231; b = 8'd73;  #10 
a = 8'd231; b = 8'd74;  #10 
a = 8'd231; b = 8'd75;  #10 
a = 8'd231; b = 8'd76;  #10 
a = 8'd231; b = 8'd77;  #10 
a = 8'd231; b = 8'd78;  #10 
a = 8'd231; b = 8'd79;  #10 
a = 8'd231; b = 8'd80;  #10 
a = 8'd231; b = 8'd81;  #10 
a = 8'd231; b = 8'd82;  #10 
a = 8'd231; b = 8'd83;  #10 
a = 8'd231; b = 8'd84;  #10 
a = 8'd231; b = 8'd85;  #10 
a = 8'd231; b = 8'd86;  #10 
a = 8'd231; b = 8'd87;  #10 
a = 8'd231; b = 8'd88;  #10 
a = 8'd231; b = 8'd89;  #10 
a = 8'd231; b = 8'd90;  #10 
a = 8'd231; b = 8'd91;  #10 
a = 8'd231; b = 8'd92;  #10 
a = 8'd231; b = 8'd93;  #10 
a = 8'd231; b = 8'd94;  #10 
a = 8'd231; b = 8'd95;  #10 
a = 8'd231; b = 8'd96;  #10 
a = 8'd231; b = 8'd97;  #10 
a = 8'd231; b = 8'd98;  #10 
a = 8'd231; b = 8'd99;  #10 
a = 8'd231; b = 8'd100;  #10 
a = 8'd231; b = 8'd101;  #10 
a = 8'd231; b = 8'd102;  #10 
a = 8'd231; b = 8'd103;  #10 
a = 8'd231; b = 8'd104;  #10 
a = 8'd231; b = 8'd105;  #10 
a = 8'd231; b = 8'd106;  #10 
a = 8'd231; b = 8'd107;  #10 
a = 8'd231; b = 8'd108;  #10 
a = 8'd231; b = 8'd109;  #10 
a = 8'd231; b = 8'd110;  #10 
a = 8'd231; b = 8'd111;  #10 
a = 8'd231; b = 8'd112;  #10 
a = 8'd231; b = 8'd113;  #10 
a = 8'd231; b = 8'd114;  #10 
a = 8'd231; b = 8'd115;  #10 
a = 8'd231; b = 8'd116;  #10 
a = 8'd231; b = 8'd117;  #10 
a = 8'd231; b = 8'd118;  #10 
a = 8'd231; b = 8'd119;  #10 
a = 8'd231; b = 8'd120;  #10 
a = 8'd231; b = 8'd121;  #10 
a = 8'd231; b = 8'd122;  #10 
a = 8'd231; b = 8'd123;  #10 
a = 8'd231; b = 8'd124;  #10 
a = 8'd231; b = 8'd125;  #10 
a = 8'd231; b = 8'd126;  #10 
a = 8'd231; b = 8'd127;  #10 
a = 8'd231; b = 8'd128;  #10 
a = 8'd231; b = 8'd129;  #10 
a = 8'd231; b = 8'd130;  #10 
a = 8'd231; b = 8'd131;  #10 
a = 8'd231; b = 8'd132;  #10 
a = 8'd231; b = 8'd133;  #10 
a = 8'd231; b = 8'd134;  #10 
a = 8'd231; b = 8'd135;  #10 
a = 8'd231; b = 8'd136;  #10 
a = 8'd231; b = 8'd137;  #10 
a = 8'd231; b = 8'd138;  #10 
a = 8'd231; b = 8'd139;  #10 
a = 8'd231; b = 8'd140;  #10 
a = 8'd231; b = 8'd141;  #10 
a = 8'd231; b = 8'd142;  #10 
a = 8'd231; b = 8'd143;  #10 
a = 8'd231; b = 8'd144;  #10 
a = 8'd231; b = 8'd145;  #10 
a = 8'd231; b = 8'd146;  #10 
a = 8'd231; b = 8'd147;  #10 
a = 8'd231; b = 8'd148;  #10 
a = 8'd231; b = 8'd149;  #10 
a = 8'd231; b = 8'd150;  #10 
a = 8'd231; b = 8'd151;  #10 
a = 8'd231; b = 8'd152;  #10 
a = 8'd231; b = 8'd153;  #10 
a = 8'd231; b = 8'd154;  #10 
a = 8'd231; b = 8'd155;  #10 
a = 8'd231; b = 8'd156;  #10 
a = 8'd231; b = 8'd157;  #10 
a = 8'd231; b = 8'd158;  #10 
a = 8'd231; b = 8'd159;  #10 
a = 8'd231; b = 8'd160;  #10 
a = 8'd231; b = 8'd161;  #10 
a = 8'd231; b = 8'd162;  #10 
a = 8'd231; b = 8'd163;  #10 
a = 8'd231; b = 8'd164;  #10 
a = 8'd231; b = 8'd165;  #10 
a = 8'd231; b = 8'd166;  #10 
a = 8'd231; b = 8'd167;  #10 
a = 8'd231; b = 8'd168;  #10 
a = 8'd231; b = 8'd169;  #10 
a = 8'd231; b = 8'd170;  #10 
a = 8'd231; b = 8'd171;  #10 
a = 8'd231; b = 8'd172;  #10 
a = 8'd231; b = 8'd173;  #10 
a = 8'd231; b = 8'd174;  #10 
a = 8'd231; b = 8'd175;  #10 
a = 8'd231; b = 8'd176;  #10 
a = 8'd231; b = 8'd177;  #10 
a = 8'd231; b = 8'd178;  #10 
a = 8'd231; b = 8'd179;  #10 
a = 8'd231; b = 8'd180;  #10 
a = 8'd231; b = 8'd181;  #10 
a = 8'd231; b = 8'd182;  #10 
a = 8'd231; b = 8'd183;  #10 
a = 8'd231; b = 8'd184;  #10 
a = 8'd231; b = 8'd185;  #10 
a = 8'd231; b = 8'd186;  #10 
a = 8'd231; b = 8'd187;  #10 
a = 8'd231; b = 8'd188;  #10 
a = 8'd231; b = 8'd189;  #10 
a = 8'd231; b = 8'd190;  #10 
a = 8'd231; b = 8'd191;  #10 
a = 8'd231; b = 8'd192;  #10 
a = 8'd231; b = 8'd193;  #10 
a = 8'd231; b = 8'd194;  #10 
a = 8'd231; b = 8'd195;  #10 
a = 8'd231; b = 8'd196;  #10 
a = 8'd231; b = 8'd197;  #10 
a = 8'd231; b = 8'd198;  #10 
a = 8'd231; b = 8'd199;  #10 
a = 8'd231; b = 8'd200;  #10 
a = 8'd231; b = 8'd201;  #10 
a = 8'd231; b = 8'd202;  #10 
a = 8'd231; b = 8'd203;  #10 
a = 8'd231; b = 8'd204;  #10 
a = 8'd231; b = 8'd205;  #10 
a = 8'd231; b = 8'd206;  #10 
a = 8'd231; b = 8'd207;  #10 
a = 8'd231; b = 8'd208;  #10 
a = 8'd231; b = 8'd209;  #10 
a = 8'd231; b = 8'd210;  #10 
a = 8'd231; b = 8'd211;  #10 
a = 8'd231; b = 8'd212;  #10 
a = 8'd231; b = 8'd213;  #10 
a = 8'd231; b = 8'd214;  #10 
a = 8'd231; b = 8'd215;  #10 
a = 8'd231; b = 8'd216;  #10 
a = 8'd231; b = 8'd217;  #10 
a = 8'd231; b = 8'd218;  #10 
a = 8'd231; b = 8'd219;  #10 
a = 8'd231; b = 8'd220;  #10 
a = 8'd231; b = 8'd221;  #10 
a = 8'd231; b = 8'd222;  #10 
a = 8'd231; b = 8'd223;  #10 
a = 8'd231; b = 8'd224;  #10 
a = 8'd231; b = 8'd225;  #10 
a = 8'd231; b = 8'd226;  #10 
a = 8'd231; b = 8'd227;  #10 
a = 8'd231; b = 8'd228;  #10 
a = 8'd231; b = 8'd229;  #10 
a = 8'd231; b = 8'd230;  #10 
a = 8'd231; b = 8'd231;  #10 
a = 8'd231; b = 8'd232;  #10 
a = 8'd231; b = 8'd233;  #10 
a = 8'd231; b = 8'd234;  #10 
a = 8'd231; b = 8'd235;  #10 
a = 8'd231; b = 8'd236;  #10 
a = 8'd231; b = 8'd237;  #10 
a = 8'd231; b = 8'd238;  #10 
a = 8'd231; b = 8'd239;  #10 
a = 8'd231; b = 8'd240;  #10 
a = 8'd231; b = 8'd241;  #10 
a = 8'd231; b = 8'd242;  #10 
a = 8'd231; b = 8'd243;  #10 
a = 8'd231; b = 8'd244;  #10 
a = 8'd231; b = 8'd245;  #10 
a = 8'd231; b = 8'd246;  #10 
a = 8'd231; b = 8'd247;  #10 
a = 8'd231; b = 8'd248;  #10 
a = 8'd231; b = 8'd249;  #10 
a = 8'd231; b = 8'd250;  #10 
a = 8'd231; b = 8'd251;  #10 
a = 8'd231; b = 8'd252;  #10 
a = 8'd231; b = 8'd253;  #10 
a = 8'd231; b = 8'd254;  #10 
a = 8'd231; b = 8'd255;  #10 
a = 8'd232; b = 8'd0;  #10 
a = 8'd232; b = 8'd1;  #10 
a = 8'd232; b = 8'd2;  #10 
a = 8'd232; b = 8'd3;  #10 
a = 8'd232; b = 8'd4;  #10 
a = 8'd232; b = 8'd5;  #10 
a = 8'd232; b = 8'd6;  #10 
a = 8'd232; b = 8'd7;  #10 
a = 8'd232; b = 8'd8;  #10 
a = 8'd232; b = 8'd9;  #10 
a = 8'd232; b = 8'd10;  #10 
a = 8'd232; b = 8'd11;  #10 
a = 8'd232; b = 8'd12;  #10 
a = 8'd232; b = 8'd13;  #10 
a = 8'd232; b = 8'd14;  #10 
a = 8'd232; b = 8'd15;  #10 
a = 8'd232; b = 8'd16;  #10 
a = 8'd232; b = 8'd17;  #10 
a = 8'd232; b = 8'd18;  #10 
a = 8'd232; b = 8'd19;  #10 
a = 8'd232; b = 8'd20;  #10 
a = 8'd232; b = 8'd21;  #10 
a = 8'd232; b = 8'd22;  #10 
a = 8'd232; b = 8'd23;  #10 
a = 8'd232; b = 8'd24;  #10 
a = 8'd232; b = 8'd25;  #10 
a = 8'd232; b = 8'd26;  #10 
a = 8'd232; b = 8'd27;  #10 
a = 8'd232; b = 8'd28;  #10 
a = 8'd232; b = 8'd29;  #10 
a = 8'd232; b = 8'd30;  #10 
a = 8'd232; b = 8'd31;  #10 
a = 8'd232; b = 8'd32;  #10 
a = 8'd232; b = 8'd33;  #10 
a = 8'd232; b = 8'd34;  #10 
a = 8'd232; b = 8'd35;  #10 
a = 8'd232; b = 8'd36;  #10 
a = 8'd232; b = 8'd37;  #10 
a = 8'd232; b = 8'd38;  #10 
a = 8'd232; b = 8'd39;  #10 
a = 8'd232; b = 8'd40;  #10 
a = 8'd232; b = 8'd41;  #10 
a = 8'd232; b = 8'd42;  #10 
a = 8'd232; b = 8'd43;  #10 
a = 8'd232; b = 8'd44;  #10 
a = 8'd232; b = 8'd45;  #10 
a = 8'd232; b = 8'd46;  #10 
a = 8'd232; b = 8'd47;  #10 
a = 8'd232; b = 8'd48;  #10 
a = 8'd232; b = 8'd49;  #10 
a = 8'd232; b = 8'd50;  #10 
a = 8'd232; b = 8'd51;  #10 
a = 8'd232; b = 8'd52;  #10 
a = 8'd232; b = 8'd53;  #10 
a = 8'd232; b = 8'd54;  #10 
a = 8'd232; b = 8'd55;  #10 
a = 8'd232; b = 8'd56;  #10 
a = 8'd232; b = 8'd57;  #10 
a = 8'd232; b = 8'd58;  #10 
a = 8'd232; b = 8'd59;  #10 
a = 8'd232; b = 8'd60;  #10 
a = 8'd232; b = 8'd61;  #10 
a = 8'd232; b = 8'd62;  #10 
a = 8'd232; b = 8'd63;  #10 
a = 8'd232; b = 8'd64;  #10 
a = 8'd232; b = 8'd65;  #10 
a = 8'd232; b = 8'd66;  #10 
a = 8'd232; b = 8'd67;  #10 
a = 8'd232; b = 8'd68;  #10 
a = 8'd232; b = 8'd69;  #10 
a = 8'd232; b = 8'd70;  #10 
a = 8'd232; b = 8'd71;  #10 
a = 8'd232; b = 8'd72;  #10 
a = 8'd232; b = 8'd73;  #10 
a = 8'd232; b = 8'd74;  #10 
a = 8'd232; b = 8'd75;  #10 
a = 8'd232; b = 8'd76;  #10 
a = 8'd232; b = 8'd77;  #10 
a = 8'd232; b = 8'd78;  #10 
a = 8'd232; b = 8'd79;  #10 
a = 8'd232; b = 8'd80;  #10 
a = 8'd232; b = 8'd81;  #10 
a = 8'd232; b = 8'd82;  #10 
a = 8'd232; b = 8'd83;  #10 
a = 8'd232; b = 8'd84;  #10 
a = 8'd232; b = 8'd85;  #10 
a = 8'd232; b = 8'd86;  #10 
a = 8'd232; b = 8'd87;  #10 
a = 8'd232; b = 8'd88;  #10 
a = 8'd232; b = 8'd89;  #10 
a = 8'd232; b = 8'd90;  #10 
a = 8'd232; b = 8'd91;  #10 
a = 8'd232; b = 8'd92;  #10 
a = 8'd232; b = 8'd93;  #10 
a = 8'd232; b = 8'd94;  #10 
a = 8'd232; b = 8'd95;  #10 
a = 8'd232; b = 8'd96;  #10 
a = 8'd232; b = 8'd97;  #10 
a = 8'd232; b = 8'd98;  #10 
a = 8'd232; b = 8'd99;  #10 
a = 8'd232; b = 8'd100;  #10 
a = 8'd232; b = 8'd101;  #10 
a = 8'd232; b = 8'd102;  #10 
a = 8'd232; b = 8'd103;  #10 
a = 8'd232; b = 8'd104;  #10 
a = 8'd232; b = 8'd105;  #10 
a = 8'd232; b = 8'd106;  #10 
a = 8'd232; b = 8'd107;  #10 
a = 8'd232; b = 8'd108;  #10 
a = 8'd232; b = 8'd109;  #10 
a = 8'd232; b = 8'd110;  #10 
a = 8'd232; b = 8'd111;  #10 
a = 8'd232; b = 8'd112;  #10 
a = 8'd232; b = 8'd113;  #10 
a = 8'd232; b = 8'd114;  #10 
a = 8'd232; b = 8'd115;  #10 
a = 8'd232; b = 8'd116;  #10 
a = 8'd232; b = 8'd117;  #10 
a = 8'd232; b = 8'd118;  #10 
a = 8'd232; b = 8'd119;  #10 
a = 8'd232; b = 8'd120;  #10 
a = 8'd232; b = 8'd121;  #10 
a = 8'd232; b = 8'd122;  #10 
a = 8'd232; b = 8'd123;  #10 
a = 8'd232; b = 8'd124;  #10 
a = 8'd232; b = 8'd125;  #10 
a = 8'd232; b = 8'd126;  #10 
a = 8'd232; b = 8'd127;  #10 
a = 8'd232; b = 8'd128;  #10 
a = 8'd232; b = 8'd129;  #10 
a = 8'd232; b = 8'd130;  #10 
a = 8'd232; b = 8'd131;  #10 
a = 8'd232; b = 8'd132;  #10 
a = 8'd232; b = 8'd133;  #10 
a = 8'd232; b = 8'd134;  #10 
a = 8'd232; b = 8'd135;  #10 
a = 8'd232; b = 8'd136;  #10 
a = 8'd232; b = 8'd137;  #10 
a = 8'd232; b = 8'd138;  #10 
a = 8'd232; b = 8'd139;  #10 
a = 8'd232; b = 8'd140;  #10 
a = 8'd232; b = 8'd141;  #10 
a = 8'd232; b = 8'd142;  #10 
a = 8'd232; b = 8'd143;  #10 
a = 8'd232; b = 8'd144;  #10 
a = 8'd232; b = 8'd145;  #10 
a = 8'd232; b = 8'd146;  #10 
a = 8'd232; b = 8'd147;  #10 
a = 8'd232; b = 8'd148;  #10 
a = 8'd232; b = 8'd149;  #10 
a = 8'd232; b = 8'd150;  #10 
a = 8'd232; b = 8'd151;  #10 
a = 8'd232; b = 8'd152;  #10 
a = 8'd232; b = 8'd153;  #10 
a = 8'd232; b = 8'd154;  #10 
a = 8'd232; b = 8'd155;  #10 
a = 8'd232; b = 8'd156;  #10 
a = 8'd232; b = 8'd157;  #10 
a = 8'd232; b = 8'd158;  #10 
a = 8'd232; b = 8'd159;  #10 
a = 8'd232; b = 8'd160;  #10 
a = 8'd232; b = 8'd161;  #10 
a = 8'd232; b = 8'd162;  #10 
a = 8'd232; b = 8'd163;  #10 
a = 8'd232; b = 8'd164;  #10 
a = 8'd232; b = 8'd165;  #10 
a = 8'd232; b = 8'd166;  #10 
a = 8'd232; b = 8'd167;  #10 
a = 8'd232; b = 8'd168;  #10 
a = 8'd232; b = 8'd169;  #10 
a = 8'd232; b = 8'd170;  #10 
a = 8'd232; b = 8'd171;  #10 
a = 8'd232; b = 8'd172;  #10 
a = 8'd232; b = 8'd173;  #10 
a = 8'd232; b = 8'd174;  #10 
a = 8'd232; b = 8'd175;  #10 
a = 8'd232; b = 8'd176;  #10 
a = 8'd232; b = 8'd177;  #10 
a = 8'd232; b = 8'd178;  #10 
a = 8'd232; b = 8'd179;  #10 
a = 8'd232; b = 8'd180;  #10 
a = 8'd232; b = 8'd181;  #10 
a = 8'd232; b = 8'd182;  #10 
a = 8'd232; b = 8'd183;  #10 
a = 8'd232; b = 8'd184;  #10 
a = 8'd232; b = 8'd185;  #10 
a = 8'd232; b = 8'd186;  #10 
a = 8'd232; b = 8'd187;  #10 
a = 8'd232; b = 8'd188;  #10 
a = 8'd232; b = 8'd189;  #10 
a = 8'd232; b = 8'd190;  #10 
a = 8'd232; b = 8'd191;  #10 
a = 8'd232; b = 8'd192;  #10 
a = 8'd232; b = 8'd193;  #10 
a = 8'd232; b = 8'd194;  #10 
a = 8'd232; b = 8'd195;  #10 
a = 8'd232; b = 8'd196;  #10 
a = 8'd232; b = 8'd197;  #10 
a = 8'd232; b = 8'd198;  #10 
a = 8'd232; b = 8'd199;  #10 
a = 8'd232; b = 8'd200;  #10 
a = 8'd232; b = 8'd201;  #10 
a = 8'd232; b = 8'd202;  #10 
a = 8'd232; b = 8'd203;  #10 
a = 8'd232; b = 8'd204;  #10 
a = 8'd232; b = 8'd205;  #10 
a = 8'd232; b = 8'd206;  #10 
a = 8'd232; b = 8'd207;  #10 
a = 8'd232; b = 8'd208;  #10 
a = 8'd232; b = 8'd209;  #10 
a = 8'd232; b = 8'd210;  #10 
a = 8'd232; b = 8'd211;  #10 
a = 8'd232; b = 8'd212;  #10 
a = 8'd232; b = 8'd213;  #10 
a = 8'd232; b = 8'd214;  #10 
a = 8'd232; b = 8'd215;  #10 
a = 8'd232; b = 8'd216;  #10 
a = 8'd232; b = 8'd217;  #10 
a = 8'd232; b = 8'd218;  #10 
a = 8'd232; b = 8'd219;  #10 
a = 8'd232; b = 8'd220;  #10 
a = 8'd232; b = 8'd221;  #10 
a = 8'd232; b = 8'd222;  #10 
a = 8'd232; b = 8'd223;  #10 
a = 8'd232; b = 8'd224;  #10 
a = 8'd232; b = 8'd225;  #10 
a = 8'd232; b = 8'd226;  #10 
a = 8'd232; b = 8'd227;  #10 
a = 8'd232; b = 8'd228;  #10 
a = 8'd232; b = 8'd229;  #10 
a = 8'd232; b = 8'd230;  #10 
a = 8'd232; b = 8'd231;  #10 
a = 8'd232; b = 8'd232;  #10 
a = 8'd232; b = 8'd233;  #10 
a = 8'd232; b = 8'd234;  #10 
a = 8'd232; b = 8'd235;  #10 
a = 8'd232; b = 8'd236;  #10 
a = 8'd232; b = 8'd237;  #10 
a = 8'd232; b = 8'd238;  #10 
a = 8'd232; b = 8'd239;  #10 
a = 8'd232; b = 8'd240;  #10 
a = 8'd232; b = 8'd241;  #10 
a = 8'd232; b = 8'd242;  #10 
a = 8'd232; b = 8'd243;  #10 
a = 8'd232; b = 8'd244;  #10 
a = 8'd232; b = 8'd245;  #10 
a = 8'd232; b = 8'd246;  #10 
a = 8'd232; b = 8'd247;  #10 
a = 8'd232; b = 8'd248;  #10 
a = 8'd232; b = 8'd249;  #10 
a = 8'd232; b = 8'd250;  #10 
a = 8'd232; b = 8'd251;  #10 
a = 8'd232; b = 8'd252;  #10 
a = 8'd232; b = 8'd253;  #10 
a = 8'd232; b = 8'd254;  #10 
a = 8'd232; b = 8'd255;  #10 
a = 8'd233; b = 8'd0;  #10 
a = 8'd233; b = 8'd1;  #10 
a = 8'd233; b = 8'd2;  #10 
a = 8'd233; b = 8'd3;  #10 
a = 8'd233; b = 8'd4;  #10 
a = 8'd233; b = 8'd5;  #10 
a = 8'd233; b = 8'd6;  #10 
a = 8'd233; b = 8'd7;  #10 
a = 8'd233; b = 8'd8;  #10 
a = 8'd233; b = 8'd9;  #10 
a = 8'd233; b = 8'd10;  #10 
a = 8'd233; b = 8'd11;  #10 
a = 8'd233; b = 8'd12;  #10 
a = 8'd233; b = 8'd13;  #10 
a = 8'd233; b = 8'd14;  #10 
a = 8'd233; b = 8'd15;  #10 
a = 8'd233; b = 8'd16;  #10 
a = 8'd233; b = 8'd17;  #10 
a = 8'd233; b = 8'd18;  #10 
a = 8'd233; b = 8'd19;  #10 
a = 8'd233; b = 8'd20;  #10 
a = 8'd233; b = 8'd21;  #10 
a = 8'd233; b = 8'd22;  #10 
a = 8'd233; b = 8'd23;  #10 
a = 8'd233; b = 8'd24;  #10 
a = 8'd233; b = 8'd25;  #10 
a = 8'd233; b = 8'd26;  #10 
a = 8'd233; b = 8'd27;  #10 
a = 8'd233; b = 8'd28;  #10 
a = 8'd233; b = 8'd29;  #10 
a = 8'd233; b = 8'd30;  #10 
a = 8'd233; b = 8'd31;  #10 
a = 8'd233; b = 8'd32;  #10 
a = 8'd233; b = 8'd33;  #10 
a = 8'd233; b = 8'd34;  #10 
a = 8'd233; b = 8'd35;  #10 
a = 8'd233; b = 8'd36;  #10 
a = 8'd233; b = 8'd37;  #10 
a = 8'd233; b = 8'd38;  #10 
a = 8'd233; b = 8'd39;  #10 
a = 8'd233; b = 8'd40;  #10 
a = 8'd233; b = 8'd41;  #10 
a = 8'd233; b = 8'd42;  #10 
a = 8'd233; b = 8'd43;  #10 
a = 8'd233; b = 8'd44;  #10 
a = 8'd233; b = 8'd45;  #10 
a = 8'd233; b = 8'd46;  #10 
a = 8'd233; b = 8'd47;  #10 
a = 8'd233; b = 8'd48;  #10 
a = 8'd233; b = 8'd49;  #10 
a = 8'd233; b = 8'd50;  #10 
a = 8'd233; b = 8'd51;  #10 
a = 8'd233; b = 8'd52;  #10 
a = 8'd233; b = 8'd53;  #10 
a = 8'd233; b = 8'd54;  #10 
a = 8'd233; b = 8'd55;  #10 
a = 8'd233; b = 8'd56;  #10 
a = 8'd233; b = 8'd57;  #10 
a = 8'd233; b = 8'd58;  #10 
a = 8'd233; b = 8'd59;  #10 
a = 8'd233; b = 8'd60;  #10 
a = 8'd233; b = 8'd61;  #10 
a = 8'd233; b = 8'd62;  #10 
a = 8'd233; b = 8'd63;  #10 
a = 8'd233; b = 8'd64;  #10 
a = 8'd233; b = 8'd65;  #10 
a = 8'd233; b = 8'd66;  #10 
a = 8'd233; b = 8'd67;  #10 
a = 8'd233; b = 8'd68;  #10 
a = 8'd233; b = 8'd69;  #10 
a = 8'd233; b = 8'd70;  #10 
a = 8'd233; b = 8'd71;  #10 
a = 8'd233; b = 8'd72;  #10 
a = 8'd233; b = 8'd73;  #10 
a = 8'd233; b = 8'd74;  #10 
a = 8'd233; b = 8'd75;  #10 
a = 8'd233; b = 8'd76;  #10 
a = 8'd233; b = 8'd77;  #10 
a = 8'd233; b = 8'd78;  #10 
a = 8'd233; b = 8'd79;  #10 
a = 8'd233; b = 8'd80;  #10 
a = 8'd233; b = 8'd81;  #10 
a = 8'd233; b = 8'd82;  #10 
a = 8'd233; b = 8'd83;  #10 
a = 8'd233; b = 8'd84;  #10 
a = 8'd233; b = 8'd85;  #10 
a = 8'd233; b = 8'd86;  #10 
a = 8'd233; b = 8'd87;  #10 
a = 8'd233; b = 8'd88;  #10 
a = 8'd233; b = 8'd89;  #10 
a = 8'd233; b = 8'd90;  #10 
a = 8'd233; b = 8'd91;  #10 
a = 8'd233; b = 8'd92;  #10 
a = 8'd233; b = 8'd93;  #10 
a = 8'd233; b = 8'd94;  #10 
a = 8'd233; b = 8'd95;  #10 
a = 8'd233; b = 8'd96;  #10 
a = 8'd233; b = 8'd97;  #10 
a = 8'd233; b = 8'd98;  #10 
a = 8'd233; b = 8'd99;  #10 
a = 8'd233; b = 8'd100;  #10 
a = 8'd233; b = 8'd101;  #10 
a = 8'd233; b = 8'd102;  #10 
a = 8'd233; b = 8'd103;  #10 
a = 8'd233; b = 8'd104;  #10 
a = 8'd233; b = 8'd105;  #10 
a = 8'd233; b = 8'd106;  #10 
a = 8'd233; b = 8'd107;  #10 
a = 8'd233; b = 8'd108;  #10 
a = 8'd233; b = 8'd109;  #10 
a = 8'd233; b = 8'd110;  #10 
a = 8'd233; b = 8'd111;  #10 
a = 8'd233; b = 8'd112;  #10 
a = 8'd233; b = 8'd113;  #10 
a = 8'd233; b = 8'd114;  #10 
a = 8'd233; b = 8'd115;  #10 
a = 8'd233; b = 8'd116;  #10 
a = 8'd233; b = 8'd117;  #10 
a = 8'd233; b = 8'd118;  #10 
a = 8'd233; b = 8'd119;  #10 
a = 8'd233; b = 8'd120;  #10 
a = 8'd233; b = 8'd121;  #10 
a = 8'd233; b = 8'd122;  #10 
a = 8'd233; b = 8'd123;  #10 
a = 8'd233; b = 8'd124;  #10 
a = 8'd233; b = 8'd125;  #10 
a = 8'd233; b = 8'd126;  #10 
a = 8'd233; b = 8'd127;  #10 
a = 8'd233; b = 8'd128;  #10 
a = 8'd233; b = 8'd129;  #10 
a = 8'd233; b = 8'd130;  #10 
a = 8'd233; b = 8'd131;  #10 
a = 8'd233; b = 8'd132;  #10 
a = 8'd233; b = 8'd133;  #10 
a = 8'd233; b = 8'd134;  #10 
a = 8'd233; b = 8'd135;  #10 
a = 8'd233; b = 8'd136;  #10 
a = 8'd233; b = 8'd137;  #10 
a = 8'd233; b = 8'd138;  #10 
a = 8'd233; b = 8'd139;  #10 
a = 8'd233; b = 8'd140;  #10 
a = 8'd233; b = 8'd141;  #10 
a = 8'd233; b = 8'd142;  #10 
a = 8'd233; b = 8'd143;  #10 
a = 8'd233; b = 8'd144;  #10 
a = 8'd233; b = 8'd145;  #10 
a = 8'd233; b = 8'd146;  #10 
a = 8'd233; b = 8'd147;  #10 
a = 8'd233; b = 8'd148;  #10 
a = 8'd233; b = 8'd149;  #10 
a = 8'd233; b = 8'd150;  #10 
a = 8'd233; b = 8'd151;  #10 
a = 8'd233; b = 8'd152;  #10 
a = 8'd233; b = 8'd153;  #10 
a = 8'd233; b = 8'd154;  #10 
a = 8'd233; b = 8'd155;  #10 
a = 8'd233; b = 8'd156;  #10 
a = 8'd233; b = 8'd157;  #10 
a = 8'd233; b = 8'd158;  #10 
a = 8'd233; b = 8'd159;  #10 
a = 8'd233; b = 8'd160;  #10 
a = 8'd233; b = 8'd161;  #10 
a = 8'd233; b = 8'd162;  #10 
a = 8'd233; b = 8'd163;  #10 
a = 8'd233; b = 8'd164;  #10 
a = 8'd233; b = 8'd165;  #10 
a = 8'd233; b = 8'd166;  #10 
a = 8'd233; b = 8'd167;  #10 
a = 8'd233; b = 8'd168;  #10 
a = 8'd233; b = 8'd169;  #10 
a = 8'd233; b = 8'd170;  #10 
a = 8'd233; b = 8'd171;  #10 
a = 8'd233; b = 8'd172;  #10 
a = 8'd233; b = 8'd173;  #10 
a = 8'd233; b = 8'd174;  #10 
a = 8'd233; b = 8'd175;  #10 
a = 8'd233; b = 8'd176;  #10 
a = 8'd233; b = 8'd177;  #10 
a = 8'd233; b = 8'd178;  #10 
a = 8'd233; b = 8'd179;  #10 
a = 8'd233; b = 8'd180;  #10 
a = 8'd233; b = 8'd181;  #10 
a = 8'd233; b = 8'd182;  #10 
a = 8'd233; b = 8'd183;  #10 
a = 8'd233; b = 8'd184;  #10 
a = 8'd233; b = 8'd185;  #10 
a = 8'd233; b = 8'd186;  #10 
a = 8'd233; b = 8'd187;  #10 
a = 8'd233; b = 8'd188;  #10 
a = 8'd233; b = 8'd189;  #10 
a = 8'd233; b = 8'd190;  #10 
a = 8'd233; b = 8'd191;  #10 
a = 8'd233; b = 8'd192;  #10 
a = 8'd233; b = 8'd193;  #10 
a = 8'd233; b = 8'd194;  #10 
a = 8'd233; b = 8'd195;  #10 
a = 8'd233; b = 8'd196;  #10 
a = 8'd233; b = 8'd197;  #10 
a = 8'd233; b = 8'd198;  #10 
a = 8'd233; b = 8'd199;  #10 
a = 8'd233; b = 8'd200;  #10 
a = 8'd233; b = 8'd201;  #10 
a = 8'd233; b = 8'd202;  #10 
a = 8'd233; b = 8'd203;  #10 
a = 8'd233; b = 8'd204;  #10 
a = 8'd233; b = 8'd205;  #10 
a = 8'd233; b = 8'd206;  #10 
a = 8'd233; b = 8'd207;  #10 
a = 8'd233; b = 8'd208;  #10 
a = 8'd233; b = 8'd209;  #10 
a = 8'd233; b = 8'd210;  #10 
a = 8'd233; b = 8'd211;  #10 
a = 8'd233; b = 8'd212;  #10 
a = 8'd233; b = 8'd213;  #10 
a = 8'd233; b = 8'd214;  #10 
a = 8'd233; b = 8'd215;  #10 
a = 8'd233; b = 8'd216;  #10 
a = 8'd233; b = 8'd217;  #10 
a = 8'd233; b = 8'd218;  #10 
a = 8'd233; b = 8'd219;  #10 
a = 8'd233; b = 8'd220;  #10 
a = 8'd233; b = 8'd221;  #10 
a = 8'd233; b = 8'd222;  #10 
a = 8'd233; b = 8'd223;  #10 
a = 8'd233; b = 8'd224;  #10 
a = 8'd233; b = 8'd225;  #10 
a = 8'd233; b = 8'd226;  #10 
a = 8'd233; b = 8'd227;  #10 
a = 8'd233; b = 8'd228;  #10 
a = 8'd233; b = 8'd229;  #10 
a = 8'd233; b = 8'd230;  #10 
a = 8'd233; b = 8'd231;  #10 
a = 8'd233; b = 8'd232;  #10 
a = 8'd233; b = 8'd233;  #10 
a = 8'd233; b = 8'd234;  #10 
a = 8'd233; b = 8'd235;  #10 
a = 8'd233; b = 8'd236;  #10 
a = 8'd233; b = 8'd237;  #10 
a = 8'd233; b = 8'd238;  #10 
a = 8'd233; b = 8'd239;  #10 
a = 8'd233; b = 8'd240;  #10 
a = 8'd233; b = 8'd241;  #10 
a = 8'd233; b = 8'd242;  #10 
a = 8'd233; b = 8'd243;  #10 
a = 8'd233; b = 8'd244;  #10 
a = 8'd233; b = 8'd245;  #10 
a = 8'd233; b = 8'd246;  #10 
a = 8'd233; b = 8'd247;  #10 
a = 8'd233; b = 8'd248;  #10 
a = 8'd233; b = 8'd249;  #10 
a = 8'd233; b = 8'd250;  #10 
a = 8'd233; b = 8'd251;  #10 
a = 8'd233; b = 8'd252;  #10 
a = 8'd233; b = 8'd253;  #10 
a = 8'd233; b = 8'd254;  #10 
a = 8'd233; b = 8'd255;  #10 
a = 8'd234; b = 8'd0;  #10 
a = 8'd234; b = 8'd1;  #10 
a = 8'd234; b = 8'd2;  #10 
a = 8'd234; b = 8'd3;  #10 
a = 8'd234; b = 8'd4;  #10 
a = 8'd234; b = 8'd5;  #10 
a = 8'd234; b = 8'd6;  #10 
a = 8'd234; b = 8'd7;  #10 
a = 8'd234; b = 8'd8;  #10 
a = 8'd234; b = 8'd9;  #10 
a = 8'd234; b = 8'd10;  #10 
a = 8'd234; b = 8'd11;  #10 
a = 8'd234; b = 8'd12;  #10 
a = 8'd234; b = 8'd13;  #10 
a = 8'd234; b = 8'd14;  #10 
a = 8'd234; b = 8'd15;  #10 
a = 8'd234; b = 8'd16;  #10 
a = 8'd234; b = 8'd17;  #10 
a = 8'd234; b = 8'd18;  #10 
a = 8'd234; b = 8'd19;  #10 
a = 8'd234; b = 8'd20;  #10 
a = 8'd234; b = 8'd21;  #10 
a = 8'd234; b = 8'd22;  #10 
a = 8'd234; b = 8'd23;  #10 
a = 8'd234; b = 8'd24;  #10 
a = 8'd234; b = 8'd25;  #10 
a = 8'd234; b = 8'd26;  #10 
a = 8'd234; b = 8'd27;  #10 
a = 8'd234; b = 8'd28;  #10 
a = 8'd234; b = 8'd29;  #10 
a = 8'd234; b = 8'd30;  #10 
a = 8'd234; b = 8'd31;  #10 
a = 8'd234; b = 8'd32;  #10 
a = 8'd234; b = 8'd33;  #10 
a = 8'd234; b = 8'd34;  #10 
a = 8'd234; b = 8'd35;  #10 
a = 8'd234; b = 8'd36;  #10 
a = 8'd234; b = 8'd37;  #10 
a = 8'd234; b = 8'd38;  #10 
a = 8'd234; b = 8'd39;  #10 
a = 8'd234; b = 8'd40;  #10 
a = 8'd234; b = 8'd41;  #10 
a = 8'd234; b = 8'd42;  #10 
a = 8'd234; b = 8'd43;  #10 
a = 8'd234; b = 8'd44;  #10 
a = 8'd234; b = 8'd45;  #10 
a = 8'd234; b = 8'd46;  #10 
a = 8'd234; b = 8'd47;  #10 
a = 8'd234; b = 8'd48;  #10 
a = 8'd234; b = 8'd49;  #10 
a = 8'd234; b = 8'd50;  #10 
a = 8'd234; b = 8'd51;  #10 
a = 8'd234; b = 8'd52;  #10 
a = 8'd234; b = 8'd53;  #10 
a = 8'd234; b = 8'd54;  #10 
a = 8'd234; b = 8'd55;  #10 
a = 8'd234; b = 8'd56;  #10 
a = 8'd234; b = 8'd57;  #10 
a = 8'd234; b = 8'd58;  #10 
a = 8'd234; b = 8'd59;  #10 
a = 8'd234; b = 8'd60;  #10 
a = 8'd234; b = 8'd61;  #10 
a = 8'd234; b = 8'd62;  #10 
a = 8'd234; b = 8'd63;  #10 
a = 8'd234; b = 8'd64;  #10 
a = 8'd234; b = 8'd65;  #10 
a = 8'd234; b = 8'd66;  #10 
a = 8'd234; b = 8'd67;  #10 
a = 8'd234; b = 8'd68;  #10 
a = 8'd234; b = 8'd69;  #10 
a = 8'd234; b = 8'd70;  #10 
a = 8'd234; b = 8'd71;  #10 
a = 8'd234; b = 8'd72;  #10 
a = 8'd234; b = 8'd73;  #10 
a = 8'd234; b = 8'd74;  #10 
a = 8'd234; b = 8'd75;  #10 
a = 8'd234; b = 8'd76;  #10 
a = 8'd234; b = 8'd77;  #10 
a = 8'd234; b = 8'd78;  #10 
a = 8'd234; b = 8'd79;  #10 
a = 8'd234; b = 8'd80;  #10 
a = 8'd234; b = 8'd81;  #10 
a = 8'd234; b = 8'd82;  #10 
a = 8'd234; b = 8'd83;  #10 
a = 8'd234; b = 8'd84;  #10 
a = 8'd234; b = 8'd85;  #10 
a = 8'd234; b = 8'd86;  #10 
a = 8'd234; b = 8'd87;  #10 
a = 8'd234; b = 8'd88;  #10 
a = 8'd234; b = 8'd89;  #10 
a = 8'd234; b = 8'd90;  #10 
a = 8'd234; b = 8'd91;  #10 
a = 8'd234; b = 8'd92;  #10 
a = 8'd234; b = 8'd93;  #10 
a = 8'd234; b = 8'd94;  #10 
a = 8'd234; b = 8'd95;  #10 
a = 8'd234; b = 8'd96;  #10 
a = 8'd234; b = 8'd97;  #10 
a = 8'd234; b = 8'd98;  #10 
a = 8'd234; b = 8'd99;  #10 
a = 8'd234; b = 8'd100;  #10 
a = 8'd234; b = 8'd101;  #10 
a = 8'd234; b = 8'd102;  #10 
a = 8'd234; b = 8'd103;  #10 
a = 8'd234; b = 8'd104;  #10 
a = 8'd234; b = 8'd105;  #10 
a = 8'd234; b = 8'd106;  #10 
a = 8'd234; b = 8'd107;  #10 
a = 8'd234; b = 8'd108;  #10 
a = 8'd234; b = 8'd109;  #10 
a = 8'd234; b = 8'd110;  #10 
a = 8'd234; b = 8'd111;  #10 
a = 8'd234; b = 8'd112;  #10 
a = 8'd234; b = 8'd113;  #10 
a = 8'd234; b = 8'd114;  #10 
a = 8'd234; b = 8'd115;  #10 
a = 8'd234; b = 8'd116;  #10 
a = 8'd234; b = 8'd117;  #10 
a = 8'd234; b = 8'd118;  #10 
a = 8'd234; b = 8'd119;  #10 
a = 8'd234; b = 8'd120;  #10 
a = 8'd234; b = 8'd121;  #10 
a = 8'd234; b = 8'd122;  #10 
a = 8'd234; b = 8'd123;  #10 
a = 8'd234; b = 8'd124;  #10 
a = 8'd234; b = 8'd125;  #10 
a = 8'd234; b = 8'd126;  #10 
a = 8'd234; b = 8'd127;  #10 
a = 8'd234; b = 8'd128;  #10 
a = 8'd234; b = 8'd129;  #10 
a = 8'd234; b = 8'd130;  #10 
a = 8'd234; b = 8'd131;  #10 
a = 8'd234; b = 8'd132;  #10 
a = 8'd234; b = 8'd133;  #10 
a = 8'd234; b = 8'd134;  #10 
a = 8'd234; b = 8'd135;  #10 
a = 8'd234; b = 8'd136;  #10 
a = 8'd234; b = 8'd137;  #10 
a = 8'd234; b = 8'd138;  #10 
a = 8'd234; b = 8'd139;  #10 
a = 8'd234; b = 8'd140;  #10 
a = 8'd234; b = 8'd141;  #10 
a = 8'd234; b = 8'd142;  #10 
a = 8'd234; b = 8'd143;  #10 
a = 8'd234; b = 8'd144;  #10 
a = 8'd234; b = 8'd145;  #10 
a = 8'd234; b = 8'd146;  #10 
a = 8'd234; b = 8'd147;  #10 
a = 8'd234; b = 8'd148;  #10 
a = 8'd234; b = 8'd149;  #10 
a = 8'd234; b = 8'd150;  #10 
a = 8'd234; b = 8'd151;  #10 
a = 8'd234; b = 8'd152;  #10 
a = 8'd234; b = 8'd153;  #10 
a = 8'd234; b = 8'd154;  #10 
a = 8'd234; b = 8'd155;  #10 
a = 8'd234; b = 8'd156;  #10 
a = 8'd234; b = 8'd157;  #10 
a = 8'd234; b = 8'd158;  #10 
a = 8'd234; b = 8'd159;  #10 
a = 8'd234; b = 8'd160;  #10 
a = 8'd234; b = 8'd161;  #10 
a = 8'd234; b = 8'd162;  #10 
a = 8'd234; b = 8'd163;  #10 
a = 8'd234; b = 8'd164;  #10 
a = 8'd234; b = 8'd165;  #10 
a = 8'd234; b = 8'd166;  #10 
a = 8'd234; b = 8'd167;  #10 
a = 8'd234; b = 8'd168;  #10 
a = 8'd234; b = 8'd169;  #10 
a = 8'd234; b = 8'd170;  #10 
a = 8'd234; b = 8'd171;  #10 
a = 8'd234; b = 8'd172;  #10 
a = 8'd234; b = 8'd173;  #10 
a = 8'd234; b = 8'd174;  #10 
a = 8'd234; b = 8'd175;  #10 
a = 8'd234; b = 8'd176;  #10 
a = 8'd234; b = 8'd177;  #10 
a = 8'd234; b = 8'd178;  #10 
a = 8'd234; b = 8'd179;  #10 
a = 8'd234; b = 8'd180;  #10 
a = 8'd234; b = 8'd181;  #10 
a = 8'd234; b = 8'd182;  #10 
a = 8'd234; b = 8'd183;  #10 
a = 8'd234; b = 8'd184;  #10 
a = 8'd234; b = 8'd185;  #10 
a = 8'd234; b = 8'd186;  #10 
a = 8'd234; b = 8'd187;  #10 
a = 8'd234; b = 8'd188;  #10 
a = 8'd234; b = 8'd189;  #10 
a = 8'd234; b = 8'd190;  #10 
a = 8'd234; b = 8'd191;  #10 
a = 8'd234; b = 8'd192;  #10 
a = 8'd234; b = 8'd193;  #10 
a = 8'd234; b = 8'd194;  #10 
a = 8'd234; b = 8'd195;  #10 
a = 8'd234; b = 8'd196;  #10 
a = 8'd234; b = 8'd197;  #10 
a = 8'd234; b = 8'd198;  #10 
a = 8'd234; b = 8'd199;  #10 
a = 8'd234; b = 8'd200;  #10 
a = 8'd234; b = 8'd201;  #10 
a = 8'd234; b = 8'd202;  #10 
a = 8'd234; b = 8'd203;  #10 
a = 8'd234; b = 8'd204;  #10 
a = 8'd234; b = 8'd205;  #10 
a = 8'd234; b = 8'd206;  #10 
a = 8'd234; b = 8'd207;  #10 
a = 8'd234; b = 8'd208;  #10 
a = 8'd234; b = 8'd209;  #10 
a = 8'd234; b = 8'd210;  #10 
a = 8'd234; b = 8'd211;  #10 
a = 8'd234; b = 8'd212;  #10 
a = 8'd234; b = 8'd213;  #10 
a = 8'd234; b = 8'd214;  #10 
a = 8'd234; b = 8'd215;  #10 
a = 8'd234; b = 8'd216;  #10 
a = 8'd234; b = 8'd217;  #10 
a = 8'd234; b = 8'd218;  #10 
a = 8'd234; b = 8'd219;  #10 
a = 8'd234; b = 8'd220;  #10 
a = 8'd234; b = 8'd221;  #10 
a = 8'd234; b = 8'd222;  #10 
a = 8'd234; b = 8'd223;  #10 
a = 8'd234; b = 8'd224;  #10 
a = 8'd234; b = 8'd225;  #10 
a = 8'd234; b = 8'd226;  #10 
a = 8'd234; b = 8'd227;  #10 
a = 8'd234; b = 8'd228;  #10 
a = 8'd234; b = 8'd229;  #10 
a = 8'd234; b = 8'd230;  #10 
a = 8'd234; b = 8'd231;  #10 
a = 8'd234; b = 8'd232;  #10 
a = 8'd234; b = 8'd233;  #10 
a = 8'd234; b = 8'd234;  #10 
a = 8'd234; b = 8'd235;  #10 
a = 8'd234; b = 8'd236;  #10 
a = 8'd234; b = 8'd237;  #10 
a = 8'd234; b = 8'd238;  #10 
a = 8'd234; b = 8'd239;  #10 
a = 8'd234; b = 8'd240;  #10 
a = 8'd234; b = 8'd241;  #10 
a = 8'd234; b = 8'd242;  #10 
a = 8'd234; b = 8'd243;  #10 
a = 8'd234; b = 8'd244;  #10 
a = 8'd234; b = 8'd245;  #10 
a = 8'd234; b = 8'd246;  #10 
a = 8'd234; b = 8'd247;  #10 
a = 8'd234; b = 8'd248;  #10 
a = 8'd234; b = 8'd249;  #10 
a = 8'd234; b = 8'd250;  #10 
a = 8'd234; b = 8'd251;  #10 
a = 8'd234; b = 8'd252;  #10 
a = 8'd234; b = 8'd253;  #10 
a = 8'd234; b = 8'd254;  #10 
a = 8'd234; b = 8'd255;  #10 
a = 8'd235; b = 8'd0;  #10 
a = 8'd235; b = 8'd1;  #10 
a = 8'd235; b = 8'd2;  #10 
a = 8'd235; b = 8'd3;  #10 
a = 8'd235; b = 8'd4;  #10 
a = 8'd235; b = 8'd5;  #10 
a = 8'd235; b = 8'd6;  #10 
a = 8'd235; b = 8'd7;  #10 
a = 8'd235; b = 8'd8;  #10 
a = 8'd235; b = 8'd9;  #10 
a = 8'd235; b = 8'd10;  #10 
a = 8'd235; b = 8'd11;  #10 
a = 8'd235; b = 8'd12;  #10 
a = 8'd235; b = 8'd13;  #10 
a = 8'd235; b = 8'd14;  #10 
a = 8'd235; b = 8'd15;  #10 
a = 8'd235; b = 8'd16;  #10 
a = 8'd235; b = 8'd17;  #10 
a = 8'd235; b = 8'd18;  #10 
a = 8'd235; b = 8'd19;  #10 
a = 8'd235; b = 8'd20;  #10 
a = 8'd235; b = 8'd21;  #10 
a = 8'd235; b = 8'd22;  #10 
a = 8'd235; b = 8'd23;  #10 
a = 8'd235; b = 8'd24;  #10 
a = 8'd235; b = 8'd25;  #10 
a = 8'd235; b = 8'd26;  #10 
a = 8'd235; b = 8'd27;  #10 
a = 8'd235; b = 8'd28;  #10 
a = 8'd235; b = 8'd29;  #10 
a = 8'd235; b = 8'd30;  #10 
a = 8'd235; b = 8'd31;  #10 
a = 8'd235; b = 8'd32;  #10 
a = 8'd235; b = 8'd33;  #10 
a = 8'd235; b = 8'd34;  #10 
a = 8'd235; b = 8'd35;  #10 
a = 8'd235; b = 8'd36;  #10 
a = 8'd235; b = 8'd37;  #10 
a = 8'd235; b = 8'd38;  #10 
a = 8'd235; b = 8'd39;  #10 
a = 8'd235; b = 8'd40;  #10 
a = 8'd235; b = 8'd41;  #10 
a = 8'd235; b = 8'd42;  #10 
a = 8'd235; b = 8'd43;  #10 
a = 8'd235; b = 8'd44;  #10 
a = 8'd235; b = 8'd45;  #10 
a = 8'd235; b = 8'd46;  #10 
a = 8'd235; b = 8'd47;  #10 
a = 8'd235; b = 8'd48;  #10 
a = 8'd235; b = 8'd49;  #10 
a = 8'd235; b = 8'd50;  #10 
a = 8'd235; b = 8'd51;  #10 
a = 8'd235; b = 8'd52;  #10 
a = 8'd235; b = 8'd53;  #10 
a = 8'd235; b = 8'd54;  #10 
a = 8'd235; b = 8'd55;  #10 
a = 8'd235; b = 8'd56;  #10 
a = 8'd235; b = 8'd57;  #10 
a = 8'd235; b = 8'd58;  #10 
a = 8'd235; b = 8'd59;  #10 
a = 8'd235; b = 8'd60;  #10 
a = 8'd235; b = 8'd61;  #10 
a = 8'd235; b = 8'd62;  #10 
a = 8'd235; b = 8'd63;  #10 
a = 8'd235; b = 8'd64;  #10 
a = 8'd235; b = 8'd65;  #10 
a = 8'd235; b = 8'd66;  #10 
a = 8'd235; b = 8'd67;  #10 
a = 8'd235; b = 8'd68;  #10 
a = 8'd235; b = 8'd69;  #10 
a = 8'd235; b = 8'd70;  #10 
a = 8'd235; b = 8'd71;  #10 
a = 8'd235; b = 8'd72;  #10 
a = 8'd235; b = 8'd73;  #10 
a = 8'd235; b = 8'd74;  #10 
a = 8'd235; b = 8'd75;  #10 
a = 8'd235; b = 8'd76;  #10 
a = 8'd235; b = 8'd77;  #10 
a = 8'd235; b = 8'd78;  #10 
a = 8'd235; b = 8'd79;  #10 
a = 8'd235; b = 8'd80;  #10 
a = 8'd235; b = 8'd81;  #10 
a = 8'd235; b = 8'd82;  #10 
a = 8'd235; b = 8'd83;  #10 
a = 8'd235; b = 8'd84;  #10 
a = 8'd235; b = 8'd85;  #10 
a = 8'd235; b = 8'd86;  #10 
a = 8'd235; b = 8'd87;  #10 
a = 8'd235; b = 8'd88;  #10 
a = 8'd235; b = 8'd89;  #10 
a = 8'd235; b = 8'd90;  #10 
a = 8'd235; b = 8'd91;  #10 
a = 8'd235; b = 8'd92;  #10 
a = 8'd235; b = 8'd93;  #10 
a = 8'd235; b = 8'd94;  #10 
a = 8'd235; b = 8'd95;  #10 
a = 8'd235; b = 8'd96;  #10 
a = 8'd235; b = 8'd97;  #10 
a = 8'd235; b = 8'd98;  #10 
a = 8'd235; b = 8'd99;  #10 
a = 8'd235; b = 8'd100;  #10 
a = 8'd235; b = 8'd101;  #10 
a = 8'd235; b = 8'd102;  #10 
a = 8'd235; b = 8'd103;  #10 
a = 8'd235; b = 8'd104;  #10 
a = 8'd235; b = 8'd105;  #10 
a = 8'd235; b = 8'd106;  #10 
a = 8'd235; b = 8'd107;  #10 
a = 8'd235; b = 8'd108;  #10 
a = 8'd235; b = 8'd109;  #10 
a = 8'd235; b = 8'd110;  #10 
a = 8'd235; b = 8'd111;  #10 
a = 8'd235; b = 8'd112;  #10 
a = 8'd235; b = 8'd113;  #10 
a = 8'd235; b = 8'd114;  #10 
a = 8'd235; b = 8'd115;  #10 
a = 8'd235; b = 8'd116;  #10 
a = 8'd235; b = 8'd117;  #10 
a = 8'd235; b = 8'd118;  #10 
a = 8'd235; b = 8'd119;  #10 
a = 8'd235; b = 8'd120;  #10 
a = 8'd235; b = 8'd121;  #10 
a = 8'd235; b = 8'd122;  #10 
a = 8'd235; b = 8'd123;  #10 
a = 8'd235; b = 8'd124;  #10 
a = 8'd235; b = 8'd125;  #10 
a = 8'd235; b = 8'd126;  #10 
a = 8'd235; b = 8'd127;  #10 
a = 8'd235; b = 8'd128;  #10 
a = 8'd235; b = 8'd129;  #10 
a = 8'd235; b = 8'd130;  #10 
a = 8'd235; b = 8'd131;  #10 
a = 8'd235; b = 8'd132;  #10 
a = 8'd235; b = 8'd133;  #10 
a = 8'd235; b = 8'd134;  #10 
a = 8'd235; b = 8'd135;  #10 
a = 8'd235; b = 8'd136;  #10 
a = 8'd235; b = 8'd137;  #10 
a = 8'd235; b = 8'd138;  #10 
a = 8'd235; b = 8'd139;  #10 
a = 8'd235; b = 8'd140;  #10 
a = 8'd235; b = 8'd141;  #10 
a = 8'd235; b = 8'd142;  #10 
a = 8'd235; b = 8'd143;  #10 
a = 8'd235; b = 8'd144;  #10 
a = 8'd235; b = 8'd145;  #10 
a = 8'd235; b = 8'd146;  #10 
a = 8'd235; b = 8'd147;  #10 
a = 8'd235; b = 8'd148;  #10 
a = 8'd235; b = 8'd149;  #10 
a = 8'd235; b = 8'd150;  #10 
a = 8'd235; b = 8'd151;  #10 
a = 8'd235; b = 8'd152;  #10 
a = 8'd235; b = 8'd153;  #10 
a = 8'd235; b = 8'd154;  #10 
a = 8'd235; b = 8'd155;  #10 
a = 8'd235; b = 8'd156;  #10 
a = 8'd235; b = 8'd157;  #10 
a = 8'd235; b = 8'd158;  #10 
a = 8'd235; b = 8'd159;  #10 
a = 8'd235; b = 8'd160;  #10 
a = 8'd235; b = 8'd161;  #10 
a = 8'd235; b = 8'd162;  #10 
a = 8'd235; b = 8'd163;  #10 
a = 8'd235; b = 8'd164;  #10 
a = 8'd235; b = 8'd165;  #10 
a = 8'd235; b = 8'd166;  #10 
a = 8'd235; b = 8'd167;  #10 
a = 8'd235; b = 8'd168;  #10 
a = 8'd235; b = 8'd169;  #10 
a = 8'd235; b = 8'd170;  #10 
a = 8'd235; b = 8'd171;  #10 
a = 8'd235; b = 8'd172;  #10 
a = 8'd235; b = 8'd173;  #10 
a = 8'd235; b = 8'd174;  #10 
a = 8'd235; b = 8'd175;  #10 
a = 8'd235; b = 8'd176;  #10 
a = 8'd235; b = 8'd177;  #10 
a = 8'd235; b = 8'd178;  #10 
a = 8'd235; b = 8'd179;  #10 
a = 8'd235; b = 8'd180;  #10 
a = 8'd235; b = 8'd181;  #10 
a = 8'd235; b = 8'd182;  #10 
a = 8'd235; b = 8'd183;  #10 
a = 8'd235; b = 8'd184;  #10 
a = 8'd235; b = 8'd185;  #10 
a = 8'd235; b = 8'd186;  #10 
a = 8'd235; b = 8'd187;  #10 
a = 8'd235; b = 8'd188;  #10 
a = 8'd235; b = 8'd189;  #10 
a = 8'd235; b = 8'd190;  #10 
a = 8'd235; b = 8'd191;  #10 
a = 8'd235; b = 8'd192;  #10 
a = 8'd235; b = 8'd193;  #10 
a = 8'd235; b = 8'd194;  #10 
a = 8'd235; b = 8'd195;  #10 
a = 8'd235; b = 8'd196;  #10 
a = 8'd235; b = 8'd197;  #10 
a = 8'd235; b = 8'd198;  #10 
a = 8'd235; b = 8'd199;  #10 
a = 8'd235; b = 8'd200;  #10 
a = 8'd235; b = 8'd201;  #10 
a = 8'd235; b = 8'd202;  #10 
a = 8'd235; b = 8'd203;  #10 
a = 8'd235; b = 8'd204;  #10 
a = 8'd235; b = 8'd205;  #10 
a = 8'd235; b = 8'd206;  #10 
a = 8'd235; b = 8'd207;  #10 
a = 8'd235; b = 8'd208;  #10 
a = 8'd235; b = 8'd209;  #10 
a = 8'd235; b = 8'd210;  #10 
a = 8'd235; b = 8'd211;  #10 
a = 8'd235; b = 8'd212;  #10 
a = 8'd235; b = 8'd213;  #10 
a = 8'd235; b = 8'd214;  #10 
a = 8'd235; b = 8'd215;  #10 
a = 8'd235; b = 8'd216;  #10 
a = 8'd235; b = 8'd217;  #10 
a = 8'd235; b = 8'd218;  #10 
a = 8'd235; b = 8'd219;  #10 
a = 8'd235; b = 8'd220;  #10 
a = 8'd235; b = 8'd221;  #10 
a = 8'd235; b = 8'd222;  #10 
a = 8'd235; b = 8'd223;  #10 
a = 8'd235; b = 8'd224;  #10 
a = 8'd235; b = 8'd225;  #10 
a = 8'd235; b = 8'd226;  #10 
a = 8'd235; b = 8'd227;  #10 
a = 8'd235; b = 8'd228;  #10 
a = 8'd235; b = 8'd229;  #10 
a = 8'd235; b = 8'd230;  #10 
a = 8'd235; b = 8'd231;  #10 
a = 8'd235; b = 8'd232;  #10 
a = 8'd235; b = 8'd233;  #10 
a = 8'd235; b = 8'd234;  #10 
a = 8'd235; b = 8'd235;  #10 
a = 8'd235; b = 8'd236;  #10 
a = 8'd235; b = 8'd237;  #10 
a = 8'd235; b = 8'd238;  #10 
a = 8'd235; b = 8'd239;  #10 
a = 8'd235; b = 8'd240;  #10 
a = 8'd235; b = 8'd241;  #10 
a = 8'd235; b = 8'd242;  #10 
a = 8'd235; b = 8'd243;  #10 
a = 8'd235; b = 8'd244;  #10 
a = 8'd235; b = 8'd245;  #10 
a = 8'd235; b = 8'd246;  #10 
a = 8'd235; b = 8'd247;  #10 
a = 8'd235; b = 8'd248;  #10 
a = 8'd235; b = 8'd249;  #10 
a = 8'd235; b = 8'd250;  #10 
a = 8'd235; b = 8'd251;  #10 
a = 8'd235; b = 8'd252;  #10 
a = 8'd235; b = 8'd253;  #10 
a = 8'd235; b = 8'd254;  #10 
a = 8'd235; b = 8'd255;  #10 
a = 8'd236; b = 8'd0;  #10 
a = 8'd236; b = 8'd1;  #10 
a = 8'd236; b = 8'd2;  #10 
a = 8'd236; b = 8'd3;  #10 
a = 8'd236; b = 8'd4;  #10 
a = 8'd236; b = 8'd5;  #10 
a = 8'd236; b = 8'd6;  #10 
a = 8'd236; b = 8'd7;  #10 
a = 8'd236; b = 8'd8;  #10 
a = 8'd236; b = 8'd9;  #10 
a = 8'd236; b = 8'd10;  #10 
a = 8'd236; b = 8'd11;  #10 
a = 8'd236; b = 8'd12;  #10 
a = 8'd236; b = 8'd13;  #10 
a = 8'd236; b = 8'd14;  #10 
a = 8'd236; b = 8'd15;  #10 
a = 8'd236; b = 8'd16;  #10 
a = 8'd236; b = 8'd17;  #10 
a = 8'd236; b = 8'd18;  #10 
a = 8'd236; b = 8'd19;  #10 
a = 8'd236; b = 8'd20;  #10 
a = 8'd236; b = 8'd21;  #10 
a = 8'd236; b = 8'd22;  #10 
a = 8'd236; b = 8'd23;  #10 
a = 8'd236; b = 8'd24;  #10 
a = 8'd236; b = 8'd25;  #10 
a = 8'd236; b = 8'd26;  #10 
a = 8'd236; b = 8'd27;  #10 
a = 8'd236; b = 8'd28;  #10 
a = 8'd236; b = 8'd29;  #10 
a = 8'd236; b = 8'd30;  #10 
a = 8'd236; b = 8'd31;  #10 
a = 8'd236; b = 8'd32;  #10 
a = 8'd236; b = 8'd33;  #10 
a = 8'd236; b = 8'd34;  #10 
a = 8'd236; b = 8'd35;  #10 
a = 8'd236; b = 8'd36;  #10 
a = 8'd236; b = 8'd37;  #10 
a = 8'd236; b = 8'd38;  #10 
a = 8'd236; b = 8'd39;  #10 
a = 8'd236; b = 8'd40;  #10 
a = 8'd236; b = 8'd41;  #10 
a = 8'd236; b = 8'd42;  #10 
a = 8'd236; b = 8'd43;  #10 
a = 8'd236; b = 8'd44;  #10 
a = 8'd236; b = 8'd45;  #10 
a = 8'd236; b = 8'd46;  #10 
a = 8'd236; b = 8'd47;  #10 
a = 8'd236; b = 8'd48;  #10 
a = 8'd236; b = 8'd49;  #10 
a = 8'd236; b = 8'd50;  #10 
a = 8'd236; b = 8'd51;  #10 
a = 8'd236; b = 8'd52;  #10 
a = 8'd236; b = 8'd53;  #10 
a = 8'd236; b = 8'd54;  #10 
a = 8'd236; b = 8'd55;  #10 
a = 8'd236; b = 8'd56;  #10 
a = 8'd236; b = 8'd57;  #10 
a = 8'd236; b = 8'd58;  #10 
a = 8'd236; b = 8'd59;  #10 
a = 8'd236; b = 8'd60;  #10 
a = 8'd236; b = 8'd61;  #10 
a = 8'd236; b = 8'd62;  #10 
a = 8'd236; b = 8'd63;  #10 
a = 8'd236; b = 8'd64;  #10 
a = 8'd236; b = 8'd65;  #10 
a = 8'd236; b = 8'd66;  #10 
a = 8'd236; b = 8'd67;  #10 
a = 8'd236; b = 8'd68;  #10 
a = 8'd236; b = 8'd69;  #10 
a = 8'd236; b = 8'd70;  #10 
a = 8'd236; b = 8'd71;  #10 
a = 8'd236; b = 8'd72;  #10 
a = 8'd236; b = 8'd73;  #10 
a = 8'd236; b = 8'd74;  #10 
a = 8'd236; b = 8'd75;  #10 
a = 8'd236; b = 8'd76;  #10 
a = 8'd236; b = 8'd77;  #10 
a = 8'd236; b = 8'd78;  #10 
a = 8'd236; b = 8'd79;  #10 
a = 8'd236; b = 8'd80;  #10 
a = 8'd236; b = 8'd81;  #10 
a = 8'd236; b = 8'd82;  #10 
a = 8'd236; b = 8'd83;  #10 
a = 8'd236; b = 8'd84;  #10 
a = 8'd236; b = 8'd85;  #10 
a = 8'd236; b = 8'd86;  #10 
a = 8'd236; b = 8'd87;  #10 
a = 8'd236; b = 8'd88;  #10 
a = 8'd236; b = 8'd89;  #10 
a = 8'd236; b = 8'd90;  #10 
a = 8'd236; b = 8'd91;  #10 
a = 8'd236; b = 8'd92;  #10 
a = 8'd236; b = 8'd93;  #10 
a = 8'd236; b = 8'd94;  #10 
a = 8'd236; b = 8'd95;  #10 
a = 8'd236; b = 8'd96;  #10 
a = 8'd236; b = 8'd97;  #10 
a = 8'd236; b = 8'd98;  #10 
a = 8'd236; b = 8'd99;  #10 
a = 8'd236; b = 8'd100;  #10 
a = 8'd236; b = 8'd101;  #10 
a = 8'd236; b = 8'd102;  #10 
a = 8'd236; b = 8'd103;  #10 
a = 8'd236; b = 8'd104;  #10 
a = 8'd236; b = 8'd105;  #10 
a = 8'd236; b = 8'd106;  #10 
a = 8'd236; b = 8'd107;  #10 
a = 8'd236; b = 8'd108;  #10 
a = 8'd236; b = 8'd109;  #10 
a = 8'd236; b = 8'd110;  #10 
a = 8'd236; b = 8'd111;  #10 
a = 8'd236; b = 8'd112;  #10 
a = 8'd236; b = 8'd113;  #10 
a = 8'd236; b = 8'd114;  #10 
a = 8'd236; b = 8'd115;  #10 
a = 8'd236; b = 8'd116;  #10 
a = 8'd236; b = 8'd117;  #10 
a = 8'd236; b = 8'd118;  #10 
a = 8'd236; b = 8'd119;  #10 
a = 8'd236; b = 8'd120;  #10 
a = 8'd236; b = 8'd121;  #10 
a = 8'd236; b = 8'd122;  #10 
a = 8'd236; b = 8'd123;  #10 
a = 8'd236; b = 8'd124;  #10 
a = 8'd236; b = 8'd125;  #10 
a = 8'd236; b = 8'd126;  #10 
a = 8'd236; b = 8'd127;  #10 
a = 8'd236; b = 8'd128;  #10 
a = 8'd236; b = 8'd129;  #10 
a = 8'd236; b = 8'd130;  #10 
a = 8'd236; b = 8'd131;  #10 
a = 8'd236; b = 8'd132;  #10 
a = 8'd236; b = 8'd133;  #10 
a = 8'd236; b = 8'd134;  #10 
a = 8'd236; b = 8'd135;  #10 
a = 8'd236; b = 8'd136;  #10 
a = 8'd236; b = 8'd137;  #10 
a = 8'd236; b = 8'd138;  #10 
a = 8'd236; b = 8'd139;  #10 
a = 8'd236; b = 8'd140;  #10 
a = 8'd236; b = 8'd141;  #10 
a = 8'd236; b = 8'd142;  #10 
a = 8'd236; b = 8'd143;  #10 
a = 8'd236; b = 8'd144;  #10 
a = 8'd236; b = 8'd145;  #10 
a = 8'd236; b = 8'd146;  #10 
a = 8'd236; b = 8'd147;  #10 
a = 8'd236; b = 8'd148;  #10 
a = 8'd236; b = 8'd149;  #10 
a = 8'd236; b = 8'd150;  #10 
a = 8'd236; b = 8'd151;  #10 
a = 8'd236; b = 8'd152;  #10 
a = 8'd236; b = 8'd153;  #10 
a = 8'd236; b = 8'd154;  #10 
a = 8'd236; b = 8'd155;  #10 
a = 8'd236; b = 8'd156;  #10 
a = 8'd236; b = 8'd157;  #10 
a = 8'd236; b = 8'd158;  #10 
a = 8'd236; b = 8'd159;  #10 
a = 8'd236; b = 8'd160;  #10 
a = 8'd236; b = 8'd161;  #10 
a = 8'd236; b = 8'd162;  #10 
a = 8'd236; b = 8'd163;  #10 
a = 8'd236; b = 8'd164;  #10 
a = 8'd236; b = 8'd165;  #10 
a = 8'd236; b = 8'd166;  #10 
a = 8'd236; b = 8'd167;  #10 
a = 8'd236; b = 8'd168;  #10 
a = 8'd236; b = 8'd169;  #10 
a = 8'd236; b = 8'd170;  #10 
a = 8'd236; b = 8'd171;  #10 
a = 8'd236; b = 8'd172;  #10 
a = 8'd236; b = 8'd173;  #10 
a = 8'd236; b = 8'd174;  #10 
a = 8'd236; b = 8'd175;  #10 
a = 8'd236; b = 8'd176;  #10 
a = 8'd236; b = 8'd177;  #10 
a = 8'd236; b = 8'd178;  #10 
a = 8'd236; b = 8'd179;  #10 
a = 8'd236; b = 8'd180;  #10 
a = 8'd236; b = 8'd181;  #10 
a = 8'd236; b = 8'd182;  #10 
a = 8'd236; b = 8'd183;  #10 
a = 8'd236; b = 8'd184;  #10 
a = 8'd236; b = 8'd185;  #10 
a = 8'd236; b = 8'd186;  #10 
a = 8'd236; b = 8'd187;  #10 
a = 8'd236; b = 8'd188;  #10 
a = 8'd236; b = 8'd189;  #10 
a = 8'd236; b = 8'd190;  #10 
a = 8'd236; b = 8'd191;  #10 
a = 8'd236; b = 8'd192;  #10 
a = 8'd236; b = 8'd193;  #10 
a = 8'd236; b = 8'd194;  #10 
a = 8'd236; b = 8'd195;  #10 
a = 8'd236; b = 8'd196;  #10 
a = 8'd236; b = 8'd197;  #10 
a = 8'd236; b = 8'd198;  #10 
a = 8'd236; b = 8'd199;  #10 
a = 8'd236; b = 8'd200;  #10 
a = 8'd236; b = 8'd201;  #10 
a = 8'd236; b = 8'd202;  #10 
a = 8'd236; b = 8'd203;  #10 
a = 8'd236; b = 8'd204;  #10 
a = 8'd236; b = 8'd205;  #10 
a = 8'd236; b = 8'd206;  #10 
a = 8'd236; b = 8'd207;  #10 
a = 8'd236; b = 8'd208;  #10 
a = 8'd236; b = 8'd209;  #10 
a = 8'd236; b = 8'd210;  #10 
a = 8'd236; b = 8'd211;  #10 
a = 8'd236; b = 8'd212;  #10 
a = 8'd236; b = 8'd213;  #10 
a = 8'd236; b = 8'd214;  #10 
a = 8'd236; b = 8'd215;  #10 
a = 8'd236; b = 8'd216;  #10 
a = 8'd236; b = 8'd217;  #10 
a = 8'd236; b = 8'd218;  #10 
a = 8'd236; b = 8'd219;  #10 
a = 8'd236; b = 8'd220;  #10 
a = 8'd236; b = 8'd221;  #10 
a = 8'd236; b = 8'd222;  #10 
a = 8'd236; b = 8'd223;  #10 
a = 8'd236; b = 8'd224;  #10 
a = 8'd236; b = 8'd225;  #10 
a = 8'd236; b = 8'd226;  #10 
a = 8'd236; b = 8'd227;  #10 
a = 8'd236; b = 8'd228;  #10 
a = 8'd236; b = 8'd229;  #10 
a = 8'd236; b = 8'd230;  #10 
a = 8'd236; b = 8'd231;  #10 
a = 8'd236; b = 8'd232;  #10 
a = 8'd236; b = 8'd233;  #10 
a = 8'd236; b = 8'd234;  #10 
a = 8'd236; b = 8'd235;  #10 
a = 8'd236; b = 8'd236;  #10 
a = 8'd236; b = 8'd237;  #10 
a = 8'd236; b = 8'd238;  #10 
a = 8'd236; b = 8'd239;  #10 
a = 8'd236; b = 8'd240;  #10 
a = 8'd236; b = 8'd241;  #10 
a = 8'd236; b = 8'd242;  #10 
a = 8'd236; b = 8'd243;  #10 
a = 8'd236; b = 8'd244;  #10 
a = 8'd236; b = 8'd245;  #10 
a = 8'd236; b = 8'd246;  #10 
a = 8'd236; b = 8'd247;  #10 
a = 8'd236; b = 8'd248;  #10 
a = 8'd236; b = 8'd249;  #10 
a = 8'd236; b = 8'd250;  #10 
a = 8'd236; b = 8'd251;  #10 
a = 8'd236; b = 8'd252;  #10 
a = 8'd236; b = 8'd253;  #10 
a = 8'd236; b = 8'd254;  #10 
a = 8'd236; b = 8'd255;  #10 
a = 8'd237; b = 8'd0;  #10 
a = 8'd237; b = 8'd1;  #10 
a = 8'd237; b = 8'd2;  #10 
a = 8'd237; b = 8'd3;  #10 
a = 8'd237; b = 8'd4;  #10 
a = 8'd237; b = 8'd5;  #10 
a = 8'd237; b = 8'd6;  #10 
a = 8'd237; b = 8'd7;  #10 
a = 8'd237; b = 8'd8;  #10 
a = 8'd237; b = 8'd9;  #10 
a = 8'd237; b = 8'd10;  #10 
a = 8'd237; b = 8'd11;  #10 
a = 8'd237; b = 8'd12;  #10 
a = 8'd237; b = 8'd13;  #10 
a = 8'd237; b = 8'd14;  #10 
a = 8'd237; b = 8'd15;  #10 
a = 8'd237; b = 8'd16;  #10 
a = 8'd237; b = 8'd17;  #10 
a = 8'd237; b = 8'd18;  #10 
a = 8'd237; b = 8'd19;  #10 
a = 8'd237; b = 8'd20;  #10 
a = 8'd237; b = 8'd21;  #10 
a = 8'd237; b = 8'd22;  #10 
a = 8'd237; b = 8'd23;  #10 
a = 8'd237; b = 8'd24;  #10 
a = 8'd237; b = 8'd25;  #10 
a = 8'd237; b = 8'd26;  #10 
a = 8'd237; b = 8'd27;  #10 
a = 8'd237; b = 8'd28;  #10 
a = 8'd237; b = 8'd29;  #10 
a = 8'd237; b = 8'd30;  #10 
a = 8'd237; b = 8'd31;  #10 
a = 8'd237; b = 8'd32;  #10 
a = 8'd237; b = 8'd33;  #10 
a = 8'd237; b = 8'd34;  #10 
a = 8'd237; b = 8'd35;  #10 
a = 8'd237; b = 8'd36;  #10 
a = 8'd237; b = 8'd37;  #10 
a = 8'd237; b = 8'd38;  #10 
a = 8'd237; b = 8'd39;  #10 
a = 8'd237; b = 8'd40;  #10 
a = 8'd237; b = 8'd41;  #10 
a = 8'd237; b = 8'd42;  #10 
a = 8'd237; b = 8'd43;  #10 
a = 8'd237; b = 8'd44;  #10 
a = 8'd237; b = 8'd45;  #10 
a = 8'd237; b = 8'd46;  #10 
a = 8'd237; b = 8'd47;  #10 
a = 8'd237; b = 8'd48;  #10 
a = 8'd237; b = 8'd49;  #10 
a = 8'd237; b = 8'd50;  #10 
a = 8'd237; b = 8'd51;  #10 
a = 8'd237; b = 8'd52;  #10 
a = 8'd237; b = 8'd53;  #10 
a = 8'd237; b = 8'd54;  #10 
a = 8'd237; b = 8'd55;  #10 
a = 8'd237; b = 8'd56;  #10 
a = 8'd237; b = 8'd57;  #10 
a = 8'd237; b = 8'd58;  #10 
a = 8'd237; b = 8'd59;  #10 
a = 8'd237; b = 8'd60;  #10 
a = 8'd237; b = 8'd61;  #10 
a = 8'd237; b = 8'd62;  #10 
a = 8'd237; b = 8'd63;  #10 
a = 8'd237; b = 8'd64;  #10 
a = 8'd237; b = 8'd65;  #10 
a = 8'd237; b = 8'd66;  #10 
a = 8'd237; b = 8'd67;  #10 
a = 8'd237; b = 8'd68;  #10 
a = 8'd237; b = 8'd69;  #10 
a = 8'd237; b = 8'd70;  #10 
a = 8'd237; b = 8'd71;  #10 
a = 8'd237; b = 8'd72;  #10 
a = 8'd237; b = 8'd73;  #10 
a = 8'd237; b = 8'd74;  #10 
a = 8'd237; b = 8'd75;  #10 
a = 8'd237; b = 8'd76;  #10 
a = 8'd237; b = 8'd77;  #10 
a = 8'd237; b = 8'd78;  #10 
a = 8'd237; b = 8'd79;  #10 
a = 8'd237; b = 8'd80;  #10 
a = 8'd237; b = 8'd81;  #10 
a = 8'd237; b = 8'd82;  #10 
a = 8'd237; b = 8'd83;  #10 
a = 8'd237; b = 8'd84;  #10 
a = 8'd237; b = 8'd85;  #10 
a = 8'd237; b = 8'd86;  #10 
a = 8'd237; b = 8'd87;  #10 
a = 8'd237; b = 8'd88;  #10 
a = 8'd237; b = 8'd89;  #10 
a = 8'd237; b = 8'd90;  #10 
a = 8'd237; b = 8'd91;  #10 
a = 8'd237; b = 8'd92;  #10 
a = 8'd237; b = 8'd93;  #10 
a = 8'd237; b = 8'd94;  #10 
a = 8'd237; b = 8'd95;  #10 
a = 8'd237; b = 8'd96;  #10 
a = 8'd237; b = 8'd97;  #10 
a = 8'd237; b = 8'd98;  #10 
a = 8'd237; b = 8'd99;  #10 
a = 8'd237; b = 8'd100;  #10 
a = 8'd237; b = 8'd101;  #10 
a = 8'd237; b = 8'd102;  #10 
a = 8'd237; b = 8'd103;  #10 
a = 8'd237; b = 8'd104;  #10 
a = 8'd237; b = 8'd105;  #10 
a = 8'd237; b = 8'd106;  #10 
a = 8'd237; b = 8'd107;  #10 
a = 8'd237; b = 8'd108;  #10 
a = 8'd237; b = 8'd109;  #10 
a = 8'd237; b = 8'd110;  #10 
a = 8'd237; b = 8'd111;  #10 
a = 8'd237; b = 8'd112;  #10 
a = 8'd237; b = 8'd113;  #10 
a = 8'd237; b = 8'd114;  #10 
a = 8'd237; b = 8'd115;  #10 
a = 8'd237; b = 8'd116;  #10 
a = 8'd237; b = 8'd117;  #10 
a = 8'd237; b = 8'd118;  #10 
a = 8'd237; b = 8'd119;  #10 
a = 8'd237; b = 8'd120;  #10 
a = 8'd237; b = 8'd121;  #10 
a = 8'd237; b = 8'd122;  #10 
a = 8'd237; b = 8'd123;  #10 
a = 8'd237; b = 8'd124;  #10 
a = 8'd237; b = 8'd125;  #10 
a = 8'd237; b = 8'd126;  #10 
a = 8'd237; b = 8'd127;  #10 
a = 8'd237; b = 8'd128;  #10 
a = 8'd237; b = 8'd129;  #10 
a = 8'd237; b = 8'd130;  #10 
a = 8'd237; b = 8'd131;  #10 
a = 8'd237; b = 8'd132;  #10 
a = 8'd237; b = 8'd133;  #10 
a = 8'd237; b = 8'd134;  #10 
a = 8'd237; b = 8'd135;  #10 
a = 8'd237; b = 8'd136;  #10 
a = 8'd237; b = 8'd137;  #10 
a = 8'd237; b = 8'd138;  #10 
a = 8'd237; b = 8'd139;  #10 
a = 8'd237; b = 8'd140;  #10 
a = 8'd237; b = 8'd141;  #10 
a = 8'd237; b = 8'd142;  #10 
a = 8'd237; b = 8'd143;  #10 
a = 8'd237; b = 8'd144;  #10 
a = 8'd237; b = 8'd145;  #10 
a = 8'd237; b = 8'd146;  #10 
a = 8'd237; b = 8'd147;  #10 
a = 8'd237; b = 8'd148;  #10 
a = 8'd237; b = 8'd149;  #10 
a = 8'd237; b = 8'd150;  #10 
a = 8'd237; b = 8'd151;  #10 
a = 8'd237; b = 8'd152;  #10 
a = 8'd237; b = 8'd153;  #10 
a = 8'd237; b = 8'd154;  #10 
a = 8'd237; b = 8'd155;  #10 
a = 8'd237; b = 8'd156;  #10 
a = 8'd237; b = 8'd157;  #10 
a = 8'd237; b = 8'd158;  #10 
a = 8'd237; b = 8'd159;  #10 
a = 8'd237; b = 8'd160;  #10 
a = 8'd237; b = 8'd161;  #10 
a = 8'd237; b = 8'd162;  #10 
a = 8'd237; b = 8'd163;  #10 
a = 8'd237; b = 8'd164;  #10 
a = 8'd237; b = 8'd165;  #10 
a = 8'd237; b = 8'd166;  #10 
a = 8'd237; b = 8'd167;  #10 
a = 8'd237; b = 8'd168;  #10 
a = 8'd237; b = 8'd169;  #10 
a = 8'd237; b = 8'd170;  #10 
a = 8'd237; b = 8'd171;  #10 
a = 8'd237; b = 8'd172;  #10 
a = 8'd237; b = 8'd173;  #10 
a = 8'd237; b = 8'd174;  #10 
a = 8'd237; b = 8'd175;  #10 
a = 8'd237; b = 8'd176;  #10 
a = 8'd237; b = 8'd177;  #10 
a = 8'd237; b = 8'd178;  #10 
a = 8'd237; b = 8'd179;  #10 
a = 8'd237; b = 8'd180;  #10 
a = 8'd237; b = 8'd181;  #10 
a = 8'd237; b = 8'd182;  #10 
a = 8'd237; b = 8'd183;  #10 
a = 8'd237; b = 8'd184;  #10 
a = 8'd237; b = 8'd185;  #10 
a = 8'd237; b = 8'd186;  #10 
a = 8'd237; b = 8'd187;  #10 
a = 8'd237; b = 8'd188;  #10 
a = 8'd237; b = 8'd189;  #10 
a = 8'd237; b = 8'd190;  #10 
a = 8'd237; b = 8'd191;  #10 
a = 8'd237; b = 8'd192;  #10 
a = 8'd237; b = 8'd193;  #10 
a = 8'd237; b = 8'd194;  #10 
a = 8'd237; b = 8'd195;  #10 
a = 8'd237; b = 8'd196;  #10 
a = 8'd237; b = 8'd197;  #10 
a = 8'd237; b = 8'd198;  #10 
a = 8'd237; b = 8'd199;  #10 
a = 8'd237; b = 8'd200;  #10 
a = 8'd237; b = 8'd201;  #10 
a = 8'd237; b = 8'd202;  #10 
a = 8'd237; b = 8'd203;  #10 
a = 8'd237; b = 8'd204;  #10 
a = 8'd237; b = 8'd205;  #10 
a = 8'd237; b = 8'd206;  #10 
a = 8'd237; b = 8'd207;  #10 
a = 8'd237; b = 8'd208;  #10 
a = 8'd237; b = 8'd209;  #10 
a = 8'd237; b = 8'd210;  #10 
a = 8'd237; b = 8'd211;  #10 
a = 8'd237; b = 8'd212;  #10 
a = 8'd237; b = 8'd213;  #10 
a = 8'd237; b = 8'd214;  #10 
a = 8'd237; b = 8'd215;  #10 
a = 8'd237; b = 8'd216;  #10 
a = 8'd237; b = 8'd217;  #10 
a = 8'd237; b = 8'd218;  #10 
a = 8'd237; b = 8'd219;  #10 
a = 8'd237; b = 8'd220;  #10 
a = 8'd237; b = 8'd221;  #10 
a = 8'd237; b = 8'd222;  #10 
a = 8'd237; b = 8'd223;  #10 
a = 8'd237; b = 8'd224;  #10 
a = 8'd237; b = 8'd225;  #10 
a = 8'd237; b = 8'd226;  #10 
a = 8'd237; b = 8'd227;  #10 
a = 8'd237; b = 8'd228;  #10 
a = 8'd237; b = 8'd229;  #10 
a = 8'd237; b = 8'd230;  #10 
a = 8'd237; b = 8'd231;  #10 
a = 8'd237; b = 8'd232;  #10 
a = 8'd237; b = 8'd233;  #10 
a = 8'd237; b = 8'd234;  #10 
a = 8'd237; b = 8'd235;  #10 
a = 8'd237; b = 8'd236;  #10 
a = 8'd237; b = 8'd237;  #10 
a = 8'd237; b = 8'd238;  #10 
a = 8'd237; b = 8'd239;  #10 
a = 8'd237; b = 8'd240;  #10 
a = 8'd237; b = 8'd241;  #10 
a = 8'd237; b = 8'd242;  #10 
a = 8'd237; b = 8'd243;  #10 
a = 8'd237; b = 8'd244;  #10 
a = 8'd237; b = 8'd245;  #10 
a = 8'd237; b = 8'd246;  #10 
a = 8'd237; b = 8'd247;  #10 
a = 8'd237; b = 8'd248;  #10 
a = 8'd237; b = 8'd249;  #10 
a = 8'd237; b = 8'd250;  #10 
a = 8'd237; b = 8'd251;  #10 
a = 8'd237; b = 8'd252;  #10 
a = 8'd237; b = 8'd253;  #10 
a = 8'd237; b = 8'd254;  #10 
a = 8'd237; b = 8'd255;  #10 
a = 8'd238; b = 8'd0;  #10 
a = 8'd238; b = 8'd1;  #10 
a = 8'd238; b = 8'd2;  #10 
a = 8'd238; b = 8'd3;  #10 
a = 8'd238; b = 8'd4;  #10 
a = 8'd238; b = 8'd5;  #10 
a = 8'd238; b = 8'd6;  #10 
a = 8'd238; b = 8'd7;  #10 
a = 8'd238; b = 8'd8;  #10 
a = 8'd238; b = 8'd9;  #10 
a = 8'd238; b = 8'd10;  #10 
a = 8'd238; b = 8'd11;  #10 
a = 8'd238; b = 8'd12;  #10 
a = 8'd238; b = 8'd13;  #10 
a = 8'd238; b = 8'd14;  #10 
a = 8'd238; b = 8'd15;  #10 
a = 8'd238; b = 8'd16;  #10 
a = 8'd238; b = 8'd17;  #10 
a = 8'd238; b = 8'd18;  #10 
a = 8'd238; b = 8'd19;  #10 
a = 8'd238; b = 8'd20;  #10 
a = 8'd238; b = 8'd21;  #10 
a = 8'd238; b = 8'd22;  #10 
a = 8'd238; b = 8'd23;  #10 
a = 8'd238; b = 8'd24;  #10 
a = 8'd238; b = 8'd25;  #10 
a = 8'd238; b = 8'd26;  #10 
a = 8'd238; b = 8'd27;  #10 
a = 8'd238; b = 8'd28;  #10 
a = 8'd238; b = 8'd29;  #10 
a = 8'd238; b = 8'd30;  #10 
a = 8'd238; b = 8'd31;  #10 
a = 8'd238; b = 8'd32;  #10 
a = 8'd238; b = 8'd33;  #10 
a = 8'd238; b = 8'd34;  #10 
a = 8'd238; b = 8'd35;  #10 
a = 8'd238; b = 8'd36;  #10 
a = 8'd238; b = 8'd37;  #10 
a = 8'd238; b = 8'd38;  #10 
a = 8'd238; b = 8'd39;  #10 
a = 8'd238; b = 8'd40;  #10 
a = 8'd238; b = 8'd41;  #10 
a = 8'd238; b = 8'd42;  #10 
a = 8'd238; b = 8'd43;  #10 
a = 8'd238; b = 8'd44;  #10 
a = 8'd238; b = 8'd45;  #10 
a = 8'd238; b = 8'd46;  #10 
a = 8'd238; b = 8'd47;  #10 
a = 8'd238; b = 8'd48;  #10 
a = 8'd238; b = 8'd49;  #10 
a = 8'd238; b = 8'd50;  #10 
a = 8'd238; b = 8'd51;  #10 
a = 8'd238; b = 8'd52;  #10 
a = 8'd238; b = 8'd53;  #10 
a = 8'd238; b = 8'd54;  #10 
a = 8'd238; b = 8'd55;  #10 
a = 8'd238; b = 8'd56;  #10 
a = 8'd238; b = 8'd57;  #10 
a = 8'd238; b = 8'd58;  #10 
a = 8'd238; b = 8'd59;  #10 
a = 8'd238; b = 8'd60;  #10 
a = 8'd238; b = 8'd61;  #10 
a = 8'd238; b = 8'd62;  #10 
a = 8'd238; b = 8'd63;  #10 
a = 8'd238; b = 8'd64;  #10 
a = 8'd238; b = 8'd65;  #10 
a = 8'd238; b = 8'd66;  #10 
a = 8'd238; b = 8'd67;  #10 
a = 8'd238; b = 8'd68;  #10 
a = 8'd238; b = 8'd69;  #10 
a = 8'd238; b = 8'd70;  #10 
a = 8'd238; b = 8'd71;  #10 
a = 8'd238; b = 8'd72;  #10 
a = 8'd238; b = 8'd73;  #10 
a = 8'd238; b = 8'd74;  #10 
a = 8'd238; b = 8'd75;  #10 
a = 8'd238; b = 8'd76;  #10 
a = 8'd238; b = 8'd77;  #10 
a = 8'd238; b = 8'd78;  #10 
a = 8'd238; b = 8'd79;  #10 
a = 8'd238; b = 8'd80;  #10 
a = 8'd238; b = 8'd81;  #10 
a = 8'd238; b = 8'd82;  #10 
a = 8'd238; b = 8'd83;  #10 
a = 8'd238; b = 8'd84;  #10 
a = 8'd238; b = 8'd85;  #10 
a = 8'd238; b = 8'd86;  #10 
a = 8'd238; b = 8'd87;  #10 
a = 8'd238; b = 8'd88;  #10 
a = 8'd238; b = 8'd89;  #10 
a = 8'd238; b = 8'd90;  #10 
a = 8'd238; b = 8'd91;  #10 
a = 8'd238; b = 8'd92;  #10 
a = 8'd238; b = 8'd93;  #10 
a = 8'd238; b = 8'd94;  #10 
a = 8'd238; b = 8'd95;  #10 
a = 8'd238; b = 8'd96;  #10 
a = 8'd238; b = 8'd97;  #10 
a = 8'd238; b = 8'd98;  #10 
a = 8'd238; b = 8'd99;  #10 
a = 8'd238; b = 8'd100;  #10 
a = 8'd238; b = 8'd101;  #10 
a = 8'd238; b = 8'd102;  #10 
a = 8'd238; b = 8'd103;  #10 
a = 8'd238; b = 8'd104;  #10 
a = 8'd238; b = 8'd105;  #10 
a = 8'd238; b = 8'd106;  #10 
a = 8'd238; b = 8'd107;  #10 
a = 8'd238; b = 8'd108;  #10 
a = 8'd238; b = 8'd109;  #10 
a = 8'd238; b = 8'd110;  #10 
a = 8'd238; b = 8'd111;  #10 
a = 8'd238; b = 8'd112;  #10 
a = 8'd238; b = 8'd113;  #10 
a = 8'd238; b = 8'd114;  #10 
a = 8'd238; b = 8'd115;  #10 
a = 8'd238; b = 8'd116;  #10 
a = 8'd238; b = 8'd117;  #10 
a = 8'd238; b = 8'd118;  #10 
a = 8'd238; b = 8'd119;  #10 
a = 8'd238; b = 8'd120;  #10 
a = 8'd238; b = 8'd121;  #10 
a = 8'd238; b = 8'd122;  #10 
a = 8'd238; b = 8'd123;  #10 
a = 8'd238; b = 8'd124;  #10 
a = 8'd238; b = 8'd125;  #10 
a = 8'd238; b = 8'd126;  #10 
a = 8'd238; b = 8'd127;  #10 
a = 8'd238; b = 8'd128;  #10 
a = 8'd238; b = 8'd129;  #10 
a = 8'd238; b = 8'd130;  #10 
a = 8'd238; b = 8'd131;  #10 
a = 8'd238; b = 8'd132;  #10 
a = 8'd238; b = 8'd133;  #10 
a = 8'd238; b = 8'd134;  #10 
a = 8'd238; b = 8'd135;  #10 
a = 8'd238; b = 8'd136;  #10 
a = 8'd238; b = 8'd137;  #10 
a = 8'd238; b = 8'd138;  #10 
a = 8'd238; b = 8'd139;  #10 
a = 8'd238; b = 8'd140;  #10 
a = 8'd238; b = 8'd141;  #10 
a = 8'd238; b = 8'd142;  #10 
a = 8'd238; b = 8'd143;  #10 
a = 8'd238; b = 8'd144;  #10 
a = 8'd238; b = 8'd145;  #10 
a = 8'd238; b = 8'd146;  #10 
a = 8'd238; b = 8'd147;  #10 
a = 8'd238; b = 8'd148;  #10 
a = 8'd238; b = 8'd149;  #10 
a = 8'd238; b = 8'd150;  #10 
a = 8'd238; b = 8'd151;  #10 
a = 8'd238; b = 8'd152;  #10 
a = 8'd238; b = 8'd153;  #10 
a = 8'd238; b = 8'd154;  #10 
a = 8'd238; b = 8'd155;  #10 
a = 8'd238; b = 8'd156;  #10 
a = 8'd238; b = 8'd157;  #10 
a = 8'd238; b = 8'd158;  #10 
a = 8'd238; b = 8'd159;  #10 
a = 8'd238; b = 8'd160;  #10 
a = 8'd238; b = 8'd161;  #10 
a = 8'd238; b = 8'd162;  #10 
a = 8'd238; b = 8'd163;  #10 
a = 8'd238; b = 8'd164;  #10 
a = 8'd238; b = 8'd165;  #10 
a = 8'd238; b = 8'd166;  #10 
a = 8'd238; b = 8'd167;  #10 
a = 8'd238; b = 8'd168;  #10 
a = 8'd238; b = 8'd169;  #10 
a = 8'd238; b = 8'd170;  #10 
a = 8'd238; b = 8'd171;  #10 
a = 8'd238; b = 8'd172;  #10 
a = 8'd238; b = 8'd173;  #10 
a = 8'd238; b = 8'd174;  #10 
a = 8'd238; b = 8'd175;  #10 
a = 8'd238; b = 8'd176;  #10 
a = 8'd238; b = 8'd177;  #10 
a = 8'd238; b = 8'd178;  #10 
a = 8'd238; b = 8'd179;  #10 
a = 8'd238; b = 8'd180;  #10 
a = 8'd238; b = 8'd181;  #10 
a = 8'd238; b = 8'd182;  #10 
a = 8'd238; b = 8'd183;  #10 
a = 8'd238; b = 8'd184;  #10 
a = 8'd238; b = 8'd185;  #10 
a = 8'd238; b = 8'd186;  #10 
a = 8'd238; b = 8'd187;  #10 
a = 8'd238; b = 8'd188;  #10 
a = 8'd238; b = 8'd189;  #10 
a = 8'd238; b = 8'd190;  #10 
a = 8'd238; b = 8'd191;  #10 
a = 8'd238; b = 8'd192;  #10 
a = 8'd238; b = 8'd193;  #10 
a = 8'd238; b = 8'd194;  #10 
a = 8'd238; b = 8'd195;  #10 
a = 8'd238; b = 8'd196;  #10 
a = 8'd238; b = 8'd197;  #10 
a = 8'd238; b = 8'd198;  #10 
a = 8'd238; b = 8'd199;  #10 
a = 8'd238; b = 8'd200;  #10 
a = 8'd238; b = 8'd201;  #10 
a = 8'd238; b = 8'd202;  #10 
a = 8'd238; b = 8'd203;  #10 
a = 8'd238; b = 8'd204;  #10 
a = 8'd238; b = 8'd205;  #10 
a = 8'd238; b = 8'd206;  #10 
a = 8'd238; b = 8'd207;  #10 
a = 8'd238; b = 8'd208;  #10 
a = 8'd238; b = 8'd209;  #10 
a = 8'd238; b = 8'd210;  #10 
a = 8'd238; b = 8'd211;  #10 
a = 8'd238; b = 8'd212;  #10 
a = 8'd238; b = 8'd213;  #10 
a = 8'd238; b = 8'd214;  #10 
a = 8'd238; b = 8'd215;  #10 
a = 8'd238; b = 8'd216;  #10 
a = 8'd238; b = 8'd217;  #10 
a = 8'd238; b = 8'd218;  #10 
a = 8'd238; b = 8'd219;  #10 
a = 8'd238; b = 8'd220;  #10 
a = 8'd238; b = 8'd221;  #10 
a = 8'd238; b = 8'd222;  #10 
a = 8'd238; b = 8'd223;  #10 
a = 8'd238; b = 8'd224;  #10 
a = 8'd238; b = 8'd225;  #10 
a = 8'd238; b = 8'd226;  #10 
a = 8'd238; b = 8'd227;  #10 
a = 8'd238; b = 8'd228;  #10 
a = 8'd238; b = 8'd229;  #10 
a = 8'd238; b = 8'd230;  #10 
a = 8'd238; b = 8'd231;  #10 
a = 8'd238; b = 8'd232;  #10 
a = 8'd238; b = 8'd233;  #10 
a = 8'd238; b = 8'd234;  #10 
a = 8'd238; b = 8'd235;  #10 
a = 8'd238; b = 8'd236;  #10 
a = 8'd238; b = 8'd237;  #10 
a = 8'd238; b = 8'd238;  #10 
a = 8'd238; b = 8'd239;  #10 
a = 8'd238; b = 8'd240;  #10 
a = 8'd238; b = 8'd241;  #10 
a = 8'd238; b = 8'd242;  #10 
a = 8'd238; b = 8'd243;  #10 
a = 8'd238; b = 8'd244;  #10 
a = 8'd238; b = 8'd245;  #10 
a = 8'd238; b = 8'd246;  #10 
a = 8'd238; b = 8'd247;  #10 
a = 8'd238; b = 8'd248;  #10 
a = 8'd238; b = 8'd249;  #10 
a = 8'd238; b = 8'd250;  #10 
a = 8'd238; b = 8'd251;  #10 
a = 8'd238; b = 8'd252;  #10 
a = 8'd238; b = 8'd253;  #10 
a = 8'd238; b = 8'd254;  #10 
a = 8'd238; b = 8'd255;  #10 
a = 8'd239; b = 8'd0;  #10 
a = 8'd239; b = 8'd1;  #10 
a = 8'd239; b = 8'd2;  #10 
a = 8'd239; b = 8'd3;  #10 
a = 8'd239; b = 8'd4;  #10 
a = 8'd239; b = 8'd5;  #10 
a = 8'd239; b = 8'd6;  #10 
a = 8'd239; b = 8'd7;  #10 
a = 8'd239; b = 8'd8;  #10 
a = 8'd239; b = 8'd9;  #10 
a = 8'd239; b = 8'd10;  #10 
a = 8'd239; b = 8'd11;  #10 
a = 8'd239; b = 8'd12;  #10 
a = 8'd239; b = 8'd13;  #10 
a = 8'd239; b = 8'd14;  #10 
a = 8'd239; b = 8'd15;  #10 
a = 8'd239; b = 8'd16;  #10 
a = 8'd239; b = 8'd17;  #10 
a = 8'd239; b = 8'd18;  #10 
a = 8'd239; b = 8'd19;  #10 
a = 8'd239; b = 8'd20;  #10 
a = 8'd239; b = 8'd21;  #10 
a = 8'd239; b = 8'd22;  #10 
a = 8'd239; b = 8'd23;  #10 
a = 8'd239; b = 8'd24;  #10 
a = 8'd239; b = 8'd25;  #10 
a = 8'd239; b = 8'd26;  #10 
a = 8'd239; b = 8'd27;  #10 
a = 8'd239; b = 8'd28;  #10 
a = 8'd239; b = 8'd29;  #10 
a = 8'd239; b = 8'd30;  #10 
a = 8'd239; b = 8'd31;  #10 
a = 8'd239; b = 8'd32;  #10 
a = 8'd239; b = 8'd33;  #10 
a = 8'd239; b = 8'd34;  #10 
a = 8'd239; b = 8'd35;  #10 
a = 8'd239; b = 8'd36;  #10 
a = 8'd239; b = 8'd37;  #10 
a = 8'd239; b = 8'd38;  #10 
a = 8'd239; b = 8'd39;  #10 
a = 8'd239; b = 8'd40;  #10 
a = 8'd239; b = 8'd41;  #10 
a = 8'd239; b = 8'd42;  #10 
a = 8'd239; b = 8'd43;  #10 
a = 8'd239; b = 8'd44;  #10 
a = 8'd239; b = 8'd45;  #10 
a = 8'd239; b = 8'd46;  #10 
a = 8'd239; b = 8'd47;  #10 
a = 8'd239; b = 8'd48;  #10 
a = 8'd239; b = 8'd49;  #10 
a = 8'd239; b = 8'd50;  #10 
a = 8'd239; b = 8'd51;  #10 
a = 8'd239; b = 8'd52;  #10 
a = 8'd239; b = 8'd53;  #10 
a = 8'd239; b = 8'd54;  #10 
a = 8'd239; b = 8'd55;  #10 
a = 8'd239; b = 8'd56;  #10 
a = 8'd239; b = 8'd57;  #10 
a = 8'd239; b = 8'd58;  #10 
a = 8'd239; b = 8'd59;  #10 
a = 8'd239; b = 8'd60;  #10 
a = 8'd239; b = 8'd61;  #10 
a = 8'd239; b = 8'd62;  #10 
a = 8'd239; b = 8'd63;  #10 
a = 8'd239; b = 8'd64;  #10 
a = 8'd239; b = 8'd65;  #10 
a = 8'd239; b = 8'd66;  #10 
a = 8'd239; b = 8'd67;  #10 
a = 8'd239; b = 8'd68;  #10 
a = 8'd239; b = 8'd69;  #10 
a = 8'd239; b = 8'd70;  #10 
a = 8'd239; b = 8'd71;  #10 
a = 8'd239; b = 8'd72;  #10 
a = 8'd239; b = 8'd73;  #10 
a = 8'd239; b = 8'd74;  #10 
a = 8'd239; b = 8'd75;  #10 
a = 8'd239; b = 8'd76;  #10 
a = 8'd239; b = 8'd77;  #10 
a = 8'd239; b = 8'd78;  #10 
a = 8'd239; b = 8'd79;  #10 
a = 8'd239; b = 8'd80;  #10 
a = 8'd239; b = 8'd81;  #10 
a = 8'd239; b = 8'd82;  #10 
a = 8'd239; b = 8'd83;  #10 
a = 8'd239; b = 8'd84;  #10 
a = 8'd239; b = 8'd85;  #10 
a = 8'd239; b = 8'd86;  #10 
a = 8'd239; b = 8'd87;  #10 
a = 8'd239; b = 8'd88;  #10 
a = 8'd239; b = 8'd89;  #10 
a = 8'd239; b = 8'd90;  #10 
a = 8'd239; b = 8'd91;  #10 
a = 8'd239; b = 8'd92;  #10 
a = 8'd239; b = 8'd93;  #10 
a = 8'd239; b = 8'd94;  #10 
a = 8'd239; b = 8'd95;  #10 
a = 8'd239; b = 8'd96;  #10 
a = 8'd239; b = 8'd97;  #10 
a = 8'd239; b = 8'd98;  #10 
a = 8'd239; b = 8'd99;  #10 
a = 8'd239; b = 8'd100;  #10 
a = 8'd239; b = 8'd101;  #10 
a = 8'd239; b = 8'd102;  #10 
a = 8'd239; b = 8'd103;  #10 
a = 8'd239; b = 8'd104;  #10 
a = 8'd239; b = 8'd105;  #10 
a = 8'd239; b = 8'd106;  #10 
a = 8'd239; b = 8'd107;  #10 
a = 8'd239; b = 8'd108;  #10 
a = 8'd239; b = 8'd109;  #10 
a = 8'd239; b = 8'd110;  #10 
a = 8'd239; b = 8'd111;  #10 
a = 8'd239; b = 8'd112;  #10 
a = 8'd239; b = 8'd113;  #10 
a = 8'd239; b = 8'd114;  #10 
a = 8'd239; b = 8'd115;  #10 
a = 8'd239; b = 8'd116;  #10 
a = 8'd239; b = 8'd117;  #10 
a = 8'd239; b = 8'd118;  #10 
a = 8'd239; b = 8'd119;  #10 
a = 8'd239; b = 8'd120;  #10 
a = 8'd239; b = 8'd121;  #10 
a = 8'd239; b = 8'd122;  #10 
a = 8'd239; b = 8'd123;  #10 
a = 8'd239; b = 8'd124;  #10 
a = 8'd239; b = 8'd125;  #10 
a = 8'd239; b = 8'd126;  #10 
a = 8'd239; b = 8'd127;  #10 
a = 8'd239; b = 8'd128;  #10 
a = 8'd239; b = 8'd129;  #10 
a = 8'd239; b = 8'd130;  #10 
a = 8'd239; b = 8'd131;  #10 
a = 8'd239; b = 8'd132;  #10 
a = 8'd239; b = 8'd133;  #10 
a = 8'd239; b = 8'd134;  #10 
a = 8'd239; b = 8'd135;  #10 
a = 8'd239; b = 8'd136;  #10 
a = 8'd239; b = 8'd137;  #10 
a = 8'd239; b = 8'd138;  #10 
a = 8'd239; b = 8'd139;  #10 
a = 8'd239; b = 8'd140;  #10 
a = 8'd239; b = 8'd141;  #10 
a = 8'd239; b = 8'd142;  #10 
a = 8'd239; b = 8'd143;  #10 
a = 8'd239; b = 8'd144;  #10 
a = 8'd239; b = 8'd145;  #10 
a = 8'd239; b = 8'd146;  #10 
a = 8'd239; b = 8'd147;  #10 
a = 8'd239; b = 8'd148;  #10 
a = 8'd239; b = 8'd149;  #10 
a = 8'd239; b = 8'd150;  #10 
a = 8'd239; b = 8'd151;  #10 
a = 8'd239; b = 8'd152;  #10 
a = 8'd239; b = 8'd153;  #10 
a = 8'd239; b = 8'd154;  #10 
a = 8'd239; b = 8'd155;  #10 
a = 8'd239; b = 8'd156;  #10 
a = 8'd239; b = 8'd157;  #10 
a = 8'd239; b = 8'd158;  #10 
a = 8'd239; b = 8'd159;  #10 
a = 8'd239; b = 8'd160;  #10 
a = 8'd239; b = 8'd161;  #10 
a = 8'd239; b = 8'd162;  #10 
a = 8'd239; b = 8'd163;  #10 
a = 8'd239; b = 8'd164;  #10 
a = 8'd239; b = 8'd165;  #10 
a = 8'd239; b = 8'd166;  #10 
a = 8'd239; b = 8'd167;  #10 
a = 8'd239; b = 8'd168;  #10 
a = 8'd239; b = 8'd169;  #10 
a = 8'd239; b = 8'd170;  #10 
a = 8'd239; b = 8'd171;  #10 
a = 8'd239; b = 8'd172;  #10 
a = 8'd239; b = 8'd173;  #10 
a = 8'd239; b = 8'd174;  #10 
a = 8'd239; b = 8'd175;  #10 
a = 8'd239; b = 8'd176;  #10 
a = 8'd239; b = 8'd177;  #10 
a = 8'd239; b = 8'd178;  #10 
a = 8'd239; b = 8'd179;  #10 
a = 8'd239; b = 8'd180;  #10 
a = 8'd239; b = 8'd181;  #10 
a = 8'd239; b = 8'd182;  #10 
a = 8'd239; b = 8'd183;  #10 
a = 8'd239; b = 8'd184;  #10 
a = 8'd239; b = 8'd185;  #10 
a = 8'd239; b = 8'd186;  #10 
a = 8'd239; b = 8'd187;  #10 
a = 8'd239; b = 8'd188;  #10 
a = 8'd239; b = 8'd189;  #10 
a = 8'd239; b = 8'd190;  #10 
a = 8'd239; b = 8'd191;  #10 
a = 8'd239; b = 8'd192;  #10 
a = 8'd239; b = 8'd193;  #10 
a = 8'd239; b = 8'd194;  #10 
a = 8'd239; b = 8'd195;  #10 
a = 8'd239; b = 8'd196;  #10 
a = 8'd239; b = 8'd197;  #10 
a = 8'd239; b = 8'd198;  #10 
a = 8'd239; b = 8'd199;  #10 
a = 8'd239; b = 8'd200;  #10 
a = 8'd239; b = 8'd201;  #10 
a = 8'd239; b = 8'd202;  #10 
a = 8'd239; b = 8'd203;  #10 
a = 8'd239; b = 8'd204;  #10 
a = 8'd239; b = 8'd205;  #10 
a = 8'd239; b = 8'd206;  #10 
a = 8'd239; b = 8'd207;  #10 
a = 8'd239; b = 8'd208;  #10 
a = 8'd239; b = 8'd209;  #10 
a = 8'd239; b = 8'd210;  #10 
a = 8'd239; b = 8'd211;  #10 
a = 8'd239; b = 8'd212;  #10 
a = 8'd239; b = 8'd213;  #10 
a = 8'd239; b = 8'd214;  #10 
a = 8'd239; b = 8'd215;  #10 
a = 8'd239; b = 8'd216;  #10 
a = 8'd239; b = 8'd217;  #10 
a = 8'd239; b = 8'd218;  #10 
a = 8'd239; b = 8'd219;  #10 
a = 8'd239; b = 8'd220;  #10 
a = 8'd239; b = 8'd221;  #10 
a = 8'd239; b = 8'd222;  #10 
a = 8'd239; b = 8'd223;  #10 
a = 8'd239; b = 8'd224;  #10 
a = 8'd239; b = 8'd225;  #10 
a = 8'd239; b = 8'd226;  #10 
a = 8'd239; b = 8'd227;  #10 
a = 8'd239; b = 8'd228;  #10 
a = 8'd239; b = 8'd229;  #10 
a = 8'd239; b = 8'd230;  #10 
a = 8'd239; b = 8'd231;  #10 
a = 8'd239; b = 8'd232;  #10 
a = 8'd239; b = 8'd233;  #10 
a = 8'd239; b = 8'd234;  #10 
a = 8'd239; b = 8'd235;  #10 
a = 8'd239; b = 8'd236;  #10 
a = 8'd239; b = 8'd237;  #10 
a = 8'd239; b = 8'd238;  #10 
a = 8'd239; b = 8'd239;  #10 
a = 8'd239; b = 8'd240;  #10 
a = 8'd239; b = 8'd241;  #10 
a = 8'd239; b = 8'd242;  #10 
a = 8'd239; b = 8'd243;  #10 
a = 8'd239; b = 8'd244;  #10 
a = 8'd239; b = 8'd245;  #10 
a = 8'd239; b = 8'd246;  #10 
a = 8'd239; b = 8'd247;  #10 
a = 8'd239; b = 8'd248;  #10 
a = 8'd239; b = 8'd249;  #10 
a = 8'd239; b = 8'd250;  #10 
a = 8'd239; b = 8'd251;  #10 
a = 8'd239; b = 8'd252;  #10 
a = 8'd239; b = 8'd253;  #10 
a = 8'd239; b = 8'd254;  #10 
a = 8'd239; b = 8'd255;  #10 
a = 8'd240; b = 8'd0;  #10 
a = 8'd240; b = 8'd1;  #10 
a = 8'd240; b = 8'd2;  #10 
a = 8'd240; b = 8'd3;  #10 
a = 8'd240; b = 8'd4;  #10 
a = 8'd240; b = 8'd5;  #10 
a = 8'd240; b = 8'd6;  #10 
a = 8'd240; b = 8'd7;  #10 
a = 8'd240; b = 8'd8;  #10 
a = 8'd240; b = 8'd9;  #10 
a = 8'd240; b = 8'd10;  #10 
a = 8'd240; b = 8'd11;  #10 
a = 8'd240; b = 8'd12;  #10 
a = 8'd240; b = 8'd13;  #10 
a = 8'd240; b = 8'd14;  #10 
a = 8'd240; b = 8'd15;  #10 
a = 8'd240; b = 8'd16;  #10 
a = 8'd240; b = 8'd17;  #10 
a = 8'd240; b = 8'd18;  #10 
a = 8'd240; b = 8'd19;  #10 
a = 8'd240; b = 8'd20;  #10 
a = 8'd240; b = 8'd21;  #10 
a = 8'd240; b = 8'd22;  #10 
a = 8'd240; b = 8'd23;  #10 
a = 8'd240; b = 8'd24;  #10 
a = 8'd240; b = 8'd25;  #10 
a = 8'd240; b = 8'd26;  #10 
a = 8'd240; b = 8'd27;  #10 
a = 8'd240; b = 8'd28;  #10 
a = 8'd240; b = 8'd29;  #10 
a = 8'd240; b = 8'd30;  #10 
a = 8'd240; b = 8'd31;  #10 
a = 8'd240; b = 8'd32;  #10 
a = 8'd240; b = 8'd33;  #10 
a = 8'd240; b = 8'd34;  #10 
a = 8'd240; b = 8'd35;  #10 
a = 8'd240; b = 8'd36;  #10 
a = 8'd240; b = 8'd37;  #10 
a = 8'd240; b = 8'd38;  #10 
a = 8'd240; b = 8'd39;  #10 
a = 8'd240; b = 8'd40;  #10 
a = 8'd240; b = 8'd41;  #10 
a = 8'd240; b = 8'd42;  #10 
a = 8'd240; b = 8'd43;  #10 
a = 8'd240; b = 8'd44;  #10 
a = 8'd240; b = 8'd45;  #10 
a = 8'd240; b = 8'd46;  #10 
a = 8'd240; b = 8'd47;  #10 
a = 8'd240; b = 8'd48;  #10 
a = 8'd240; b = 8'd49;  #10 
a = 8'd240; b = 8'd50;  #10 
a = 8'd240; b = 8'd51;  #10 
a = 8'd240; b = 8'd52;  #10 
a = 8'd240; b = 8'd53;  #10 
a = 8'd240; b = 8'd54;  #10 
a = 8'd240; b = 8'd55;  #10 
a = 8'd240; b = 8'd56;  #10 
a = 8'd240; b = 8'd57;  #10 
a = 8'd240; b = 8'd58;  #10 
a = 8'd240; b = 8'd59;  #10 
a = 8'd240; b = 8'd60;  #10 
a = 8'd240; b = 8'd61;  #10 
a = 8'd240; b = 8'd62;  #10 
a = 8'd240; b = 8'd63;  #10 
a = 8'd240; b = 8'd64;  #10 
a = 8'd240; b = 8'd65;  #10 
a = 8'd240; b = 8'd66;  #10 
a = 8'd240; b = 8'd67;  #10 
a = 8'd240; b = 8'd68;  #10 
a = 8'd240; b = 8'd69;  #10 
a = 8'd240; b = 8'd70;  #10 
a = 8'd240; b = 8'd71;  #10 
a = 8'd240; b = 8'd72;  #10 
a = 8'd240; b = 8'd73;  #10 
a = 8'd240; b = 8'd74;  #10 
a = 8'd240; b = 8'd75;  #10 
a = 8'd240; b = 8'd76;  #10 
a = 8'd240; b = 8'd77;  #10 
a = 8'd240; b = 8'd78;  #10 
a = 8'd240; b = 8'd79;  #10 
a = 8'd240; b = 8'd80;  #10 
a = 8'd240; b = 8'd81;  #10 
a = 8'd240; b = 8'd82;  #10 
a = 8'd240; b = 8'd83;  #10 
a = 8'd240; b = 8'd84;  #10 
a = 8'd240; b = 8'd85;  #10 
a = 8'd240; b = 8'd86;  #10 
a = 8'd240; b = 8'd87;  #10 
a = 8'd240; b = 8'd88;  #10 
a = 8'd240; b = 8'd89;  #10 
a = 8'd240; b = 8'd90;  #10 
a = 8'd240; b = 8'd91;  #10 
a = 8'd240; b = 8'd92;  #10 
a = 8'd240; b = 8'd93;  #10 
a = 8'd240; b = 8'd94;  #10 
a = 8'd240; b = 8'd95;  #10 
a = 8'd240; b = 8'd96;  #10 
a = 8'd240; b = 8'd97;  #10 
a = 8'd240; b = 8'd98;  #10 
a = 8'd240; b = 8'd99;  #10 
a = 8'd240; b = 8'd100;  #10 
a = 8'd240; b = 8'd101;  #10 
a = 8'd240; b = 8'd102;  #10 
a = 8'd240; b = 8'd103;  #10 
a = 8'd240; b = 8'd104;  #10 
a = 8'd240; b = 8'd105;  #10 
a = 8'd240; b = 8'd106;  #10 
a = 8'd240; b = 8'd107;  #10 
a = 8'd240; b = 8'd108;  #10 
a = 8'd240; b = 8'd109;  #10 
a = 8'd240; b = 8'd110;  #10 
a = 8'd240; b = 8'd111;  #10 
a = 8'd240; b = 8'd112;  #10 
a = 8'd240; b = 8'd113;  #10 
a = 8'd240; b = 8'd114;  #10 
a = 8'd240; b = 8'd115;  #10 
a = 8'd240; b = 8'd116;  #10 
a = 8'd240; b = 8'd117;  #10 
a = 8'd240; b = 8'd118;  #10 
a = 8'd240; b = 8'd119;  #10 
a = 8'd240; b = 8'd120;  #10 
a = 8'd240; b = 8'd121;  #10 
a = 8'd240; b = 8'd122;  #10 
a = 8'd240; b = 8'd123;  #10 
a = 8'd240; b = 8'd124;  #10 
a = 8'd240; b = 8'd125;  #10 
a = 8'd240; b = 8'd126;  #10 
a = 8'd240; b = 8'd127;  #10 
a = 8'd240; b = 8'd128;  #10 
a = 8'd240; b = 8'd129;  #10 
a = 8'd240; b = 8'd130;  #10 
a = 8'd240; b = 8'd131;  #10 
a = 8'd240; b = 8'd132;  #10 
a = 8'd240; b = 8'd133;  #10 
a = 8'd240; b = 8'd134;  #10 
a = 8'd240; b = 8'd135;  #10 
a = 8'd240; b = 8'd136;  #10 
a = 8'd240; b = 8'd137;  #10 
a = 8'd240; b = 8'd138;  #10 
a = 8'd240; b = 8'd139;  #10 
a = 8'd240; b = 8'd140;  #10 
a = 8'd240; b = 8'd141;  #10 
a = 8'd240; b = 8'd142;  #10 
a = 8'd240; b = 8'd143;  #10 
a = 8'd240; b = 8'd144;  #10 
a = 8'd240; b = 8'd145;  #10 
a = 8'd240; b = 8'd146;  #10 
a = 8'd240; b = 8'd147;  #10 
a = 8'd240; b = 8'd148;  #10 
a = 8'd240; b = 8'd149;  #10 
a = 8'd240; b = 8'd150;  #10 
a = 8'd240; b = 8'd151;  #10 
a = 8'd240; b = 8'd152;  #10 
a = 8'd240; b = 8'd153;  #10 
a = 8'd240; b = 8'd154;  #10 
a = 8'd240; b = 8'd155;  #10 
a = 8'd240; b = 8'd156;  #10 
a = 8'd240; b = 8'd157;  #10 
a = 8'd240; b = 8'd158;  #10 
a = 8'd240; b = 8'd159;  #10 
a = 8'd240; b = 8'd160;  #10 
a = 8'd240; b = 8'd161;  #10 
a = 8'd240; b = 8'd162;  #10 
a = 8'd240; b = 8'd163;  #10 
a = 8'd240; b = 8'd164;  #10 
a = 8'd240; b = 8'd165;  #10 
a = 8'd240; b = 8'd166;  #10 
a = 8'd240; b = 8'd167;  #10 
a = 8'd240; b = 8'd168;  #10 
a = 8'd240; b = 8'd169;  #10 
a = 8'd240; b = 8'd170;  #10 
a = 8'd240; b = 8'd171;  #10 
a = 8'd240; b = 8'd172;  #10 
a = 8'd240; b = 8'd173;  #10 
a = 8'd240; b = 8'd174;  #10 
a = 8'd240; b = 8'd175;  #10 
a = 8'd240; b = 8'd176;  #10 
a = 8'd240; b = 8'd177;  #10 
a = 8'd240; b = 8'd178;  #10 
a = 8'd240; b = 8'd179;  #10 
a = 8'd240; b = 8'd180;  #10 
a = 8'd240; b = 8'd181;  #10 
a = 8'd240; b = 8'd182;  #10 
a = 8'd240; b = 8'd183;  #10 
a = 8'd240; b = 8'd184;  #10 
a = 8'd240; b = 8'd185;  #10 
a = 8'd240; b = 8'd186;  #10 
a = 8'd240; b = 8'd187;  #10 
a = 8'd240; b = 8'd188;  #10 
a = 8'd240; b = 8'd189;  #10 
a = 8'd240; b = 8'd190;  #10 
a = 8'd240; b = 8'd191;  #10 
a = 8'd240; b = 8'd192;  #10 
a = 8'd240; b = 8'd193;  #10 
a = 8'd240; b = 8'd194;  #10 
a = 8'd240; b = 8'd195;  #10 
a = 8'd240; b = 8'd196;  #10 
a = 8'd240; b = 8'd197;  #10 
a = 8'd240; b = 8'd198;  #10 
a = 8'd240; b = 8'd199;  #10 
a = 8'd240; b = 8'd200;  #10 
a = 8'd240; b = 8'd201;  #10 
a = 8'd240; b = 8'd202;  #10 
a = 8'd240; b = 8'd203;  #10 
a = 8'd240; b = 8'd204;  #10 
a = 8'd240; b = 8'd205;  #10 
a = 8'd240; b = 8'd206;  #10 
a = 8'd240; b = 8'd207;  #10 
a = 8'd240; b = 8'd208;  #10 
a = 8'd240; b = 8'd209;  #10 
a = 8'd240; b = 8'd210;  #10 
a = 8'd240; b = 8'd211;  #10 
a = 8'd240; b = 8'd212;  #10 
a = 8'd240; b = 8'd213;  #10 
a = 8'd240; b = 8'd214;  #10 
a = 8'd240; b = 8'd215;  #10 
a = 8'd240; b = 8'd216;  #10 
a = 8'd240; b = 8'd217;  #10 
a = 8'd240; b = 8'd218;  #10 
a = 8'd240; b = 8'd219;  #10 
a = 8'd240; b = 8'd220;  #10 
a = 8'd240; b = 8'd221;  #10 
a = 8'd240; b = 8'd222;  #10 
a = 8'd240; b = 8'd223;  #10 
a = 8'd240; b = 8'd224;  #10 
a = 8'd240; b = 8'd225;  #10 
a = 8'd240; b = 8'd226;  #10 
a = 8'd240; b = 8'd227;  #10 
a = 8'd240; b = 8'd228;  #10 
a = 8'd240; b = 8'd229;  #10 
a = 8'd240; b = 8'd230;  #10 
a = 8'd240; b = 8'd231;  #10 
a = 8'd240; b = 8'd232;  #10 
a = 8'd240; b = 8'd233;  #10 
a = 8'd240; b = 8'd234;  #10 
a = 8'd240; b = 8'd235;  #10 
a = 8'd240; b = 8'd236;  #10 
a = 8'd240; b = 8'd237;  #10 
a = 8'd240; b = 8'd238;  #10 
a = 8'd240; b = 8'd239;  #10 
a = 8'd240; b = 8'd240;  #10 
a = 8'd240; b = 8'd241;  #10 
a = 8'd240; b = 8'd242;  #10 
a = 8'd240; b = 8'd243;  #10 
a = 8'd240; b = 8'd244;  #10 
a = 8'd240; b = 8'd245;  #10 
a = 8'd240; b = 8'd246;  #10 
a = 8'd240; b = 8'd247;  #10 
a = 8'd240; b = 8'd248;  #10 
a = 8'd240; b = 8'd249;  #10 
a = 8'd240; b = 8'd250;  #10 
a = 8'd240; b = 8'd251;  #10 
a = 8'd240; b = 8'd252;  #10 
a = 8'd240; b = 8'd253;  #10 
a = 8'd240; b = 8'd254;  #10 
a = 8'd240; b = 8'd255;  #10 
a = 8'd241; b = 8'd0;  #10 
a = 8'd241; b = 8'd1;  #10 
a = 8'd241; b = 8'd2;  #10 
a = 8'd241; b = 8'd3;  #10 
a = 8'd241; b = 8'd4;  #10 
a = 8'd241; b = 8'd5;  #10 
a = 8'd241; b = 8'd6;  #10 
a = 8'd241; b = 8'd7;  #10 
a = 8'd241; b = 8'd8;  #10 
a = 8'd241; b = 8'd9;  #10 
a = 8'd241; b = 8'd10;  #10 
a = 8'd241; b = 8'd11;  #10 
a = 8'd241; b = 8'd12;  #10 
a = 8'd241; b = 8'd13;  #10 
a = 8'd241; b = 8'd14;  #10 
a = 8'd241; b = 8'd15;  #10 
a = 8'd241; b = 8'd16;  #10 
a = 8'd241; b = 8'd17;  #10 
a = 8'd241; b = 8'd18;  #10 
a = 8'd241; b = 8'd19;  #10 
a = 8'd241; b = 8'd20;  #10 
a = 8'd241; b = 8'd21;  #10 
a = 8'd241; b = 8'd22;  #10 
a = 8'd241; b = 8'd23;  #10 
a = 8'd241; b = 8'd24;  #10 
a = 8'd241; b = 8'd25;  #10 
a = 8'd241; b = 8'd26;  #10 
a = 8'd241; b = 8'd27;  #10 
a = 8'd241; b = 8'd28;  #10 
a = 8'd241; b = 8'd29;  #10 
a = 8'd241; b = 8'd30;  #10 
a = 8'd241; b = 8'd31;  #10 
a = 8'd241; b = 8'd32;  #10 
a = 8'd241; b = 8'd33;  #10 
a = 8'd241; b = 8'd34;  #10 
a = 8'd241; b = 8'd35;  #10 
a = 8'd241; b = 8'd36;  #10 
a = 8'd241; b = 8'd37;  #10 
a = 8'd241; b = 8'd38;  #10 
a = 8'd241; b = 8'd39;  #10 
a = 8'd241; b = 8'd40;  #10 
a = 8'd241; b = 8'd41;  #10 
a = 8'd241; b = 8'd42;  #10 
a = 8'd241; b = 8'd43;  #10 
a = 8'd241; b = 8'd44;  #10 
a = 8'd241; b = 8'd45;  #10 
a = 8'd241; b = 8'd46;  #10 
a = 8'd241; b = 8'd47;  #10 
a = 8'd241; b = 8'd48;  #10 
a = 8'd241; b = 8'd49;  #10 
a = 8'd241; b = 8'd50;  #10 
a = 8'd241; b = 8'd51;  #10 
a = 8'd241; b = 8'd52;  #10 
a = 8'd241; b = 8'd53;  #10 
a = 8'd241; b = 8'd54;  #10 
a = 8'd241; b = 8'd55;  #10 
a = 8'd241; b = 8'd56;  #10 
a = 8'd241; b = 8'd57;  #10 
a = 8'd241; b = 8'd58;  #10 
a = 8'd241; b = 8'd59;  #10 
a = 8'd241; b = 8'd60;  #10 
a = 8'd241; b = 8'd61;  #10 
a = 8'd241; b = 8'd62;  #10 
a = 8'd241; b = 8'd63;  #10 
a = 8'd241; b = 8'd64;  #10 
a = 8'd241; b = 8'd65;  #10 
a = 8'd241; b = 8'd66;  #10 
a = 8'd241; b = 8'd67;  #10 
a = 8'd241; b = 8'd68;  #10 
a = 8'd241; b = 8'd69;  #10 
a = 8'd241; b = 8'd70;  #10 
a = 8'd241; b = 8'd71;  #10 
a = 8'd241; b = 8'd72;  #10 
a = 8'd241; b = 8'd73;  #10 
a = 8'd241; b = 8'd74;  #10 
a = 8'd241; b = 8'd75;  #10 
a = 8'd241; b = 8'd76;  #10 
a = 8'd241; b = 8'd77;  #10 
a = 8'd241; b = 8'd78;  #10 
a = 8'd241; b = 8'd79;  #10 
a = 8'd241; b = 8'd80;  #10 
a = 8'd241; b = 8'd81;  #10 
a = 8'd241; b = 8'd82;  #10 
a = 8'd241; b = 8'd83;  #10 
a = 8'd241; b = 8'd84;  #10 
a = 8'd241; b = 8'd85;  #10 
a = 8'd241; b = 8'd86;  #10 
a = 8'd241; b = 8'd87;  #10 
a = 8'd241; b = 8'd88;  #10 
a = 8'd241; b = 8'd89;  #10 
a = 8'd241; b = 8'd90;  #10 
a = 8'd241; b = 8'd91;  #10 
a = 8'd241; b = 8'd92;  #10 
a = 8'd241; b = 8'd93;  #10 
a = 8'd241; b = 8'd94;  #10 
a = 8'd241; b = 8'd95;  #10 
a = 8'd241; b = 8'd96;  #10 
a = 8'd241; b = 8'd97;  #10 
a = 8'd241; b = 8'd98;  #10 
a = 8'd241; b = 8'd99;  #10 
a = 8'd241; b = 8'd100;  #10 
a = 8'd241; b = 8'd101;  #10 
a = 8'd241; b = 8'd102;  #10 
a = 8'd241; b = 8'd103;  #10 
a = 8'd241; b = 8'd104;  #10 
a = 8'd241; b = 8'd105;  #10 
a = 8'd241; b = 8'd106;  #10 
a = 8'd241; b = 8'd107;  #10 
a = 8'd241; b = 8'd108;  #10 
a = 8'd241; b = 8'd109;  #10 
a = 8'd241; b = 8'd110;  #10 
a = 8'd241; b = 8'd111;  #10 
a = 8'd241; b = 8'd112;  #10 
a = 8'd241; b = 8'd113;  #10 
a = 8'd241; b = 8'd114;  #10 
a = 8'd241; b = 8'd115;  #10 
a = 8'd241; b = 8'd116;  #10 
a = 8'd241; b = 8'd117;  #10 
a = 8'd241; b = 8'd118;  #10 
a = 8'd241; b = 8'd119;  #10 
a = 8'd241; b = 8'd120;  #10 
a = 8'd241; b = 8'd121;  #10 
a = 8'd241; b = 8'd122;  #10 
a = 8'd241; b = 8'd123;  #10 
a = 8'd241; b = 8'd124;  #10 
a = 8'd241; b = 8'd125;  #10 
a = 8'd241; b = 8'd126;  #10 
a = 8'd241; b = 8'd127;  #10 
a = 8'd241; b = 8'd128;  #10 
a = 8'd241; b = 8'd129;  #10 
a = 8'd241; b = 8'd130;  #10 
a = 8'd241; b = 8'd131;  #10 
a = 8'd241; b = 8'd132;  #10 
a = 8'd241; b = 8'd133;  #10 
a = 8'd241; b = 8'd134;  #10 
a = 8'd241; b = 8'd135;  #10 
a = 8'd241; b = 8'd136;  #10 
a = 8'd241; b = 8'd137;  #10 
a = 8'd241; b = 8'd138;  #10 
a = 8'd241; b = 8'd139;  #10 
a = 8'd241; b = 8'd140;  #10 
a = 8'd241; b = 8'd141;  #10 
a = 8'd241; b = 8'd142;  #10 
a = 8'd241; b = 8'd143;  #10 
a = 8'd241; b = 8'd144;  #10 
a = 8'd241; b = 8'd145;  #10 
a = 8'd241; b = 8'd146;  #10 
a = 8'd241; b = 8'd147;  #10 
a = 8'd241; b = 8'd148;  #10 
a = 8'd241; b = 8'd149;  #10 
a = 8'd241; b = 8'd150;  #10 
a = 8'd241; b = 8'd151;  #10 
a = 8'd241; b = 8'd152;  #10 
a = 8'd241; b = 8'd153;  #10 
a = 8'd241; b = 8'd154;  #10 
a = 8'd241; b = 8'd155;  #10 
a = 8'd241; b = 8'd156;  #10 
a = 8'd241; b = 8'd157;  #10 
a = 8'd241; b = 8'd158;  #10 
a = 8'd241; b = 8'd159;  #10 
a = 8'd241; b = 8'd160;  #10 
a = 8'd241; b = 8'd161;  #10 
a = 8'd241; b = 8'd162;  #10 
a = 8'd241; b = 8'd163;  #10 
a = 8'd241; b = 8'd164;  #10 
a = 8'd241; b = 8'd165;  #10 
a = 8'd241; b = 8'd166;  #10 
a = 8'd241; b = 8'd167;  #10 
a = 8'd241; b = 8'd168;  #10 
a = 8'd241; b = 8'd169;  #10 
a = 8'd241; b = 8'd170;  #10 
a = 8'd241; b = 8'd171;  #10 
a = 8'd241; b = 8'd172;  #10 
a = 8'd241; b = 8'd173;  #10 
a = 8'd241; b = 8'd174;  #10 
a = 8'd241; b = 8'd175;  #10 
a = 8'd241; b = 8'd176;  #10 
a = 8'd241; b = 8'd177;  #10 
a = 8'd241; b = 8'd178;  #10 
a = 8'd241; b = 8'd179;  #10 
a = 8'd241; b = 8'd180;  #10 
a = 8'd241; b = 8'd181;  #10 
a = 8'd241; b = 8'd182;  #10 
a = 8'd241; b = 8'd183;  #10 
a = 8'd241; b = 8'd184;  #10 
a = 8'd241; b = 8'd185;  #10 
a = 8'd241; b = 8'd186;  #10 
a = 8'd241; b = 8'd187;  #10 
a = 8'd241; b = 8'd188;  #10 
a = 8'd241; b = 8'd189;  #10 
a = 8'd241; b = 8'd190;  #10 
a = 8'd241; b = 8'd191;  #10 
a = 8'd241; b = 8'd192;  #10 
a = 8'd241; b = 8'd193;  #10 
a = 8'd241; b = 8'd194;  #10 
a = 8'd241; b = 8'd195;  #10 
a = 8'd241; b = 8'd196;  #10 
a = 8'd241; b = 8'd197;  #10 
a = 8'd241; b = 8'd198;  #10 
a = 8'd241; b = 8'd199;  #10 
a = 8'd241; b = 8'd200;  #10 
a = 8'd241; b = 8'd201;  #10 
a = 8'd241; b = 8'd202;  #10 
a = 8'd241; b = 8'd203;  #10 
a = 8'd241; b = 8'd204;  #10 
a = 8'd241; b = 8'd205;  #10 
a = 8'd241; b = 8'd206;  #10 
a = 8'd241; b = 8'd207;  #10 
a = 8'd241; b = 8'd208;  #10 
a = 8'd241; b = 8'd209;  #10 
a = 8'd241; b = 8'd210;  #10 
a = 8'd241; b = 8'd211;  #10 
a = 8'd241; b = 8'd212;  #10 
a = 8'd241; b = 8'd213;  #10 
a = 8'd241; b = 8'd214;  #10 
a = 8'd241; b = 8'd215;  #10 
a = 8'd241; b = 8'd216;  #10 
a = 8'd241; b = 8'd217;  #10 
a = 8'd241; b = 8'd218;  #10 
a = 8'd241; b = 8'd219;  #10 
a = 8'd241; b = 8'd220;  #10 
a = 8'd241; b = 8'd221;  #10 
a = 8'd241; b = 8'd222;  #10 
a = 8'd241; b = 8'd223;  #10 
a = 8'd241; b = 8'd224;  #10 
a = 8'd241; b = 8'd225;  #10 
a = 8'd241; b = 8'd226;  #10 
a = 8'd241; b = 8'd227;  #10 
a = 8'd241; b = 8'd228;  #10 
a = 8'd241; b = 8'd229;  #10 
a = 8'd241; b = 8'd230;  #10 
a = 8'd241; b = 8'd231;  #10 
a = 8'd241; b = 8'd232;  #10 
a = 8'd241; b = 8'd233;  #10 
a = 8'd241; b = 8'd234;  #10 
a = 8'd241; b = 8'd235;  #10 
a = 8'd241; b = 8'd236;  #10 
a = 8'd241; b = 8'd237;  #10 
a = 8'd241; b = 8'd238;  #10 
a = 8'd241; b = 8'd239;  #10 
a = 8'd241; b = 8'd240;  #10 
a = 8'd241; b = 8'd241;  #10 
a = 8'd241; b = 8'd242;  #10 
a = 8'd241; b = 8'd243;  #10 
a = 8'd241; b = 8'd244;  #10 
a = 8'd241; b = 8'd245;  #10 
a = 8'd241; b = 8'd246;  #10 
a = 8'd241; b = 8'd247;  #10 
a = 8'd241; b = 8'd248;  #10 
a = 8'd241; b = 8'd249;  #10 
a = 8'd241; b = 8'd250;  #10 
a = 8'd241; b = 8'd251;  #10 
a = 8'd241; b = 8'd252;  #10 
a = 8'd241; b = 8'd253;  #10 
a = 8'd241; b = 8'd254;  #10 
a = 8'd241; b = 8'd255;  #10 
a = 8'd242; b = 8'd0;  #10 
a = 8'd242; b = 8'd1;  #10 
a = 8'd242; b = 8'd2;  #10 
a = 8'd242; b = 8'd3;  #10 
a = 8'd242; b = 8'd4;  #10 
a = 8'd242; b = 8'd5;  #10 
a = 8'd242; b = 8'd6;  #10 
a = 8'd242; b = 8'd7;  #10 
a = 8'd242; b = 8'd8;  #10 
a = 8'd242; b = 8'd9;  #10 
a = 8'd242; b = 8'd10;  #10 
a = 8'd242; b = 8'd11;  #10 
a = 8'd242; b = 8'd12;  #10 
a = 8'd242; b = 8'd13;  #10 
a = 8'd242; b = 8'd14;  #10 
a = 8'd242; b = 8'd15;  #10 
a = 8'd242; b = 8'd16;  #10 
a = 8'd242; b = 8'd17;  #10 
a = 8'd242; b = 8'd18;  #10 
a = 8'd242; b = 8'd19;  #10 
a = 8'd242; b = 8'd20;  #10 
a = 8'd242; b = 8'd21;  #10 
a = 8'd242; b = 8'd22;  #10 
a = 8'd242; b = 8'd23;  #10 
a = 8'd242; b = 8'd24;  #10 
a = 8'd242; b = 8'd25;  #10 
a = 8'd242; b = 8'd26;  #10 
a = 8'd242; b = 8'd27;  #10 
a = 8'd242; b = 8'd28;  #10 
a = 8'd242; b = 8'd29;  #10 
a = 8'd242; b = 8'd30;  #10 
a = 8'd242; b = 8'd31;  #10 
a = 8'd242; b = 8'd32;  #10 
a = 8'd242; b = 8'd33;  #10 
a = 8'd242; b = 8'd34;  #10 
a = 8'd242; b = 8'd35;  #10 
a = 8'd242; b = 8'd36;  #10 
a = 8'd242; b = 8'd37;  #10 
a = 8'd242; b = 8'd38;  #10 
a = 8'd242; b = 8'd39;  #10 
a = 8'd242; b = 8'd40;  #10 
a = 8'd242; b = 8'd41;  #10 
a = 8'd242; b = 8'd42;  #10 
a = 8'd242; b = 8'd43;  #10 
a = 8'd242; b = 8'd44;  #10 
a = 8'd242; b = 8'd45;  #10 
a = 8'd242; b = 8'd46;  #10 
a = 8'd242; b = 8'd47;  #10 
a = 8'd242; b = 8'd48;  #10 
a = 8'd242; b = 8'd49;  #10 
a = 8'd242; b = 8'd50;  #10 
a = 8'd242; b = 8'd51;  #10 
a = 8'd242; b = 8'd52;  #10 
a = 8'd242; b = 8'd53;  #10 
a = 8'd242; b = 8'd54;  #10 
a = 8'd242; b = 8'd55;  #10 
a = 8'd242; b = 8'd56;  #10 
a = 8'd242; b = 8'd57;  #10 
a = 8'd242; b = 8'd58;  #10 
a = 8'd242; b = 8'd59;  #10 
a = 8'd242; b = 8'd60;  #10 
a = 8'd242; b = 8'd61;  #10 
a = 8'd242; b = 8'd62;  #10 
a = 8'd242; b = 8'd63;  #10 
a = 8'd242; b = 8'd64;  #10 
a = 8'd242; b = 8'd65;  #10 
a = 8'd242; b = 8'd66;  #10 
a = 8'd242; b = 8'd67;  #10 
a = 8'd242; b = 8'd68;  #10 
a = 8'd242; b = 8'd69;  #10 
a = 8'd242; b = 8'd70;  #10 
a = 8'd242; b = 8'd71;  #10 
a = 8'd242; b = 8'd72;  #10 
a = 8'd242; b = 8'd73;  #10 
a = 8'd242; b = 8'd74;  #10 
a = 8'd242; b = 8'd75;  #10 
a = 8'd242; b = 8'd76;  #10 
a = 8'd242; b = 8'd77;  #10 
a = 8'd242; b = 8'd78;  #10 
a = 8'd242; b = 8'd79;  #10 
a = 8'd242; b = 8'd80;  #10 
a = 8'd242; b = 8'd81;  #10 
a = 8'd242; b = 8'd82;  #10 
a = 8'd242; b = 8'd83;  #10 
a = 8'd242; b = 8'd84;  #10 
a = 8'd242; b = 8'd85;  #10 
a = 8'd242; b = 8'd86;  #10 
a = 8'd242; b = 8'd87;  #10 
a = 8'd242; b = 8'd88;  #10 
a = 8'd242; b = 8'd89;  #10 
a = 8'd242; b = 8'd90;  #10 
a = 8'd242; b = 8'd91;  #10 
a = 8'd242; b = 8'd92;  #10 
a = 8'd242; b = 8'd93;  #10 
a = 8'd242; b = 8'd94;  #10 
a = 8'd242; b = 8'd95;  #10 
a = 8'd242; b = 8'd96;  #10 
a = 8'd242; b = 8'd97;  #10 
a = 8'd242; b = 8'd98;  #10 
a = 8'd242; b = 8'd99;  #10 
a = 8'd242; b = 8'd100;  #10 
a = 8'd242; b = 8'd101;  #10 
a = 8'd242; b = 8'd102;  #10 
a = 8'd242; b = 8'd103;  #10 
a = 8'd242; b = 8'd104;  #10 
a = 8'd242; b = 8'd105;  #10 
a = 8'd242; b = 8'd106;  #10 
a = 8'd242; b = 8'd107;  #10 
a = 8'd242; b = 8'd108;  #10 
a = 8'd242; b = 8'd109;  #10 
a = 8'd242; b = 8'd110;  #10 
a = 8'd242; b = 8'd111;  #10 
a = 8'd242; b = 8'd112;  #10 
a = 8'd242; b = 8'd113;  #10 
a = 8'd242; b = 8'd114;  #10 
a = 8'd242; b = 8'd115;  #10 
a = 8'd242; b = 8'd116;  #10 
a = 8'd242; b = 8'd117;  #10 
a = 8'd242; b = 8'd118;  #10 
a = 8'd242; b = 8'd119;  #10 
a = 8'd242; b = 8'd120;  #10 
a = 8'd242; b = 8'd121;  #10 
a = 8'd242; b = 8'd122;  #10 
a = 8'd242; b = 8'd123;  #10 
a = 8'd242; b = 8'd124;  #10 
a = 8'd242; b = 8'd125;  #10 
a = 8'd242; b = 8'd126;  #10 
a = 8'd242; b = 8'd127;  #10 
a = 8'd242; b = 8'd128;  #10 
a = 8'd242; b = 8'd129;  #10 
a = 8'd242; b = 8'd130;  #10 
a = 8'd242; b = 8'd131;  #10 
a = 8'd242; b = 8'd132;  #10 
a = 8'd242; b = 8'd133;  #10 
a = 8'd242; b = 8'd134;  #10 
a = 8'd242; b = 8'd135;  #10 
a = 8'd242; b = 8'd136;  #10 
a = 8'd242; b = 8'd137;  #10 
a = 8'd242; b = 8'd138;  #10 
a = 8'd242; b = 8'd139;  #10 
a = 8'd242; b = 8'd140;  #10 
a = 8'd242; b = 8'd141;  #10 
a = 8'd242; b = 8'd142;  #10 
a = 8'd242; b = 8'd143;  #10 
a = 8'd242; b = 8'd144;  #10 
a = 8'd242; b = 8'd145;  #10 
a = 8'd242; b = 8'd146;  #10 
a = 8'd242; b = 8'd147;  #10 
a = 8'd242; b = 8'd148;  #10 
a = 8'd242; b = 8'd149;  #10 
a = 8'd242; b = 8'd150;  #10 
a = 8'd242; b = 8'd151;  #10 
a = 8'd242; b = 8'd152;  #10 
a = 8'd242; b = 8'd153;  #10 
a = 8'd242; b = 8'd154;  #10 
a = 8'd242; b = 8'd155;  #10 
a = 8'd242; b = 8'd156;  #10 
a = 8'd242; b = 8'd157;  #10 
a = 8'd242; b = 8'd158;  #10 
a = 8'd242; b = 8'd159;  #10 
a = 8'd242; b = 8'd160;  #10 
a = 8'd242; b = 8'd161;  #10 
a = 8'd242; b = 8'd162;  #10 
a = 8'd242; b = 8'd163;  #10 
a = 8'd242; b = 8'd164;  #10 
a = 8'd242; b = 8'd165;  #10 
a = 8'd242; b = 8'd166;  #10 
a = 8'd242; b = 8'd167;  #10 
a = 8'd242; b = 8'd168;  #10 
a = 8'd242; b = 8'd169;  #10 
a = 8'd242; b = 8'd170;  #10 
a = 8'd242; b = 8'd171;  #10 
a = 8'd242; b = 8'd172;  #10 
a = 8'd242; b = 8'd173;  #10 
a = 8'd242; b = 8'd174;  #10 
a = 8'd242; b = 8'd175;  #10 
a = 8'd242; b = 8'd176;  #10 
a = 8'd242; b = 8'd177;  #10 
a = 8'd242; b = 8'd178;  #10 
a = 8'd242; b = 8'd179;  #10 
a = 8'd242; b = 8'd180;  #10 
a = 8'd242; b = 8'd181;  #10 
a = 8'd242; b = 8'd182;  #10 
a = 8'd242; b = 8'd183;  #10 
a = 8'd242; b = 8'd184;  #10 
a = 8'd242; b = 8'd185;  #10 
a = 8'd242; b = 8'd186;  #10 
a = 8'd242; b = 8'd187;  #10 
a = 8'd242; b = 8'd188;  #10 
a = 8'd242; b = 8'd189;  #10 
a = 8'd242; b = 8'd190;  #10 
a = 8'd242; b = 8'd191;  #10 
a = 8'd242; b = 8'd192;  #10 
a = 8'd242; b = 8'd193;  #10 
a = 8'd242; b = 8'd194;  #10 
a = 8'd242; b = 8'd195;  #10 
a = 8'd242; b = 8'd196;  #10 
a = 8'd242; b = 8'd197;  #10 
a = 8'd242; b = 8'd198;  #10 
a = 8'd242; b = 8'd199;  #10 
a = 8'd242; b = 8'd200;  #10 
a = 8'd242; b = 8'd201;  #10 
a = 8'd242; b = 8'd202;  #10 
a = 8'd242; b = 8'd203;  #10 
a = 8'd242; b = 8'd204;  #10 
a = 8'd242; b = 8'd205;  #10 
a = 8'd242; b = 8'd206;  #10 
a = 8'd242; b = 8'd207;  #10 
a = 8'd242; b = 8'd208;  #10 
a = 8'd242; b = 8'd209;  #10 
a = 8'd242; b = 8'd210;  #10 
a = 8'd242; b = 8'd211;  #10 
a = 8'd242; b = 8'd212;  #10 
a = 8'd242; b = 8'd213;  #10 
a = 8'd242; b = 8'd214;  #10 
a = 8'd242; b = 8'd215;  #10 
a = 8'd242; b = 8'd216;  #10 
a = 8'd242; b = 8'd217;  #10 
a = 8'd242; b = 8'd218;  #10 
a = 8'd242; b = 8'd219;  #10 
a = 8'd242; b = 8'd220;  #10 
a = 8'd242; b = 8'd221;  #10 
a = 8'd242; b = 8'd222;  #10 
a = 8'd242; b = 8'd223;  #10 
a = 8'd242; b = 8'd224;  #10 
a = 8'd242; b = 8'd225;  #10 
a = 8'd242; b = 8'd226;  #10 
a = 8'd242; b = 8'd227;  #10 
a = 8'd242; b = 8'd228;  #10 
a = 8'd242; b = 8'd229;  #10 
a = 8'd242; b = 8'd230;  #10 
a = 8'd242; b = 8'd231;  #10 
a = 8'd242; b = 8'd232;  #10 
a = 8'd242; b = 8'd233;  #10 
a = 8'd242; b = 8'd234;  #10 
a = 8'd242; b = 8'd235;  #10 
a = 8'd242; b = 8'd236;  #10 
a = 8'd242; b = 8'd237;  #10 
a = 8'd242; b = 8'd238;  #10 
a = 8'd242; b = 8'd239;  #10 
a = 8'd242; b = 8'd240;  #10 
a = 8'd242; b = 8'd241;  #10 
a = 8'd242; b = 8'd242;  #10 
a = 8'd242; b = 8'd243;  #10 
a = 8'd242; b = 8'd244;  #10 
a = 8'd242; b = 8'd245;  #10 
a = 8'd242; b = 8'd246;  #10 
a = 8'd242; b = 8'd247;  #10 
a = 8'd242; b = 8'd248;  #10 
a = 8'd242; b = 8'd249;  #10 
a = 8'd242; b = 8'd250;  #10 
a = 8'd242; b = 8'd251;  #10 
a = 8'd242; b = 8'd252;  #10 
a = 8'd242; b = 8'd253;  #10 
a = 8'd242; b = 8'd254;  #10 
a = 8'd242; b = 8'd255;  #10 
a = 8'd243; b = 8'd0;  #10 
a = 8'd243; b = 8'd1;  #10 
a = 8'd243; b = 8'd2;  #10 
a = 8'd243; b = 8'd3;  #10 
a = 8'd243; b = 8'd4;  #10 
a = 8'd243; b = 8'd5;  #10 
a = 8'd243; b = 8'd6;  #10 
a = 8'd243; b = 8'd7;  #10 
a = 8'd243; b = 8'd8;  #10 
a = 8'd243; b = 8'd9;  #10 
a = 8'd243; b = 8'd10;  #10 
a = 8'd243; b = 8'd11;  #10 
a = 8'd243; b = 8'd12;  #10 
a = 8'd243; b = 8'd13;  #10 
a = 8'd243; b = 8'd14;  #10 
a = 8'd243; b = 8'd15;  #10 
a = 8'd243; b = 8'd16;  #10 
a = 8'd243; b = 8'd17;  #10 
a = 8'd243; b = 8'd18;  #10 
a = 8'd243; b = 8'd19;  #10 
a = 8'd243; b = 8'd20;  #10 
a = 8'd243; b = 8'd21;  #10 
a = 8'd243; b = 8'd22;  #10 
a = 8'd243; b = 8'd23;  #10 
a = 8'd243; b = 8'd24;  #10 
a = 8'd243; b = 8'd25;  #10 
a = 8'd243; b = 8'd26;  #10 
a = 8'd243; b = 8'd27;  #10 
a = 8'd243; b = 8'd28;  #10 
a = 8'd243; b = 8'd29;  #10 
a = 8'd243; b = 8'd30;  #10 
a = 8'd243; b = 8'd31;  #10 
a = 8'd243; b = 8'd32;  #10 
a = 8'd243; b = 8'd33;  #10 
a = 8'd243; b = 8'd34;  #10 
a = 8'd243; b = 8'd35;  #10 
a = 8'd243; b = 8'd36;  #10 
a = 8'd243; b = 8'd37;  #10 
a = 8'd243; b = 8'd38;  #10 
a = 8'd243; b = 8'd39;  #10 
a = 8'd243; b = 8'd40;  #10 
a = 8'd243; b = 8'd41;  #10 
a = 8'd243; b = 8'd42;  #10 
a = 8'd243; b = 8'd43;  #10 
a = 8'd243; b = 8'd44;  #10 
a = 8'd243; b = 8'd45;  #10 
a = 8'd243; b = 8'd46;  #10 
a = 8'd243; b = 8'd47;  #10 
a = 8'd243; b = 8'd48;  #10 
a = 8'd243; b = 8'd49;  #10 
a = 8'd243; b = 8'd50;  #10 
a = 8'd243; b = 8'd51;  #10 
a = 8'd243; b = 8'd52;  #10 
a = 8'd243; b = 8'd53;  #10 
a = 8'd243; b = 8'd54;  #10 
a = 8'd243; b = 8'd55;  #10 
a = 8'd243; b = 8'd56;  #10 
a = 8'd243; b = 8'd57;  #10 
a = 8'd243; b = 8'd58;  #10 
a = 8'd243; b = 8'd59;  #10 
a = 8'd243; b = 8'd60;  #10 
a = 8'd243; b = 8'd61;  #10 
a = 8'd243; b = 8'd62;  #10 
a = 8'd243; b = 8'd63;  #10 
a = 8'd243; b = 8'd64;  #10 
a = 8'd243; b = 8'd65;  #10 
a = 8'd243; b = 8'd66;  #10 
a = 8'd243; b = 8'd67;  #10 
a = 8'd243; b = 8'd68;  #10 
a = 8'd243; b = 8'd69;  #10 
a = 8'd243; b = 8'd70;  #10 
a = 8'd243; b = 8'd71;  #10 
a = 8'd243; b = 8'd72;  #10 
a = 8'd243; b = 8'd73;  #10 
a = 8'd243; b = 8'd74;  #10 
a = 8'd243; b = 8'd75;  #10 
a = 8'd243; b = 8'd76;  #10 
a = 8'd243; b = 8'd77;  #10 
a = 8'd243; b = 8'd78;  #10 
a = 8'd243; b = 8'd79;  #10 
a = 8'd243; b = 8'd80;  #10 
a = 8'd243; b = 8'd81;  #10 
a = 8'd243; b = 8'd82;  #10 
a = 8'd243; b = 8'd83;  #10 
a = 8'd243; b = 8'd84;  #10 
a = 8'd243; b = 8'd85;  #10 
a = 8'd243; b = 8'd86;  #10 
a = 8'd243; b = 8'd87;  #10 
a = 8'd243; b = 8'd88;  #10 
a = 8'd243; b = 8'd89;  #10 
a = 8'd243; b = 8'd90;  #10 
a = 8'd243; b = 8'd91;  #10 
a = 8'd243; b = 8'd92;  #10 
a = 8'd243; b = 8'd93;  #10 
a = 8'd243; b = 8'd94;  #10 
a = 8'd243; b = 8'd95;  #10 
a = 8'd243; b = 8'd96;  #10 
a = 8'd243; b = 8'd97;  #10 
a = 8'd243; b = 8'd98;  #10 
a = 8'd243; b = 8'd99;  #10 
a = 8'd243; b = 8'd100;  #10 
a = 8'd243; b = 8'd101;  #10 
a = 8'd243; b = 8'd102;  #10 
a = 8'd243; b = 8'd103;  #10 
a = 8'd243; b = 8'd104;  #10 
a = 8'd243; b = 8'd105;  #10 
a = 8'd243; b = 8'd106;  #10 
a = 8'd243; b = 8'd107;  #10 
a = 8'd243; b = 8'd108;  #10 
a = 8'd243; b = 8'd109;  #10 
a = 8'd243; b = 8'd110;  #10 
a = 8'd243; b = 8'd111;  #10 
a = 8'd243; b = 8'd112;  #10 
a = 8'd243; b = 8'd113;  #10 
a = 8'd243; b = 8'd114;  #10 
a = 8'd243; b = 8'd115;  #10 
a = 8'd243; b = 8'd116;  #10 
a = 8'd243; b = 8'd117;  #10 
a = 8'd243; b = 8'd118;  #10 
a = 8'd243; b = 8'd119;  #10 
a = 8'd243; b = 8'd120;  #10 
a = 8'd243; b = 8'd121;  #10 
a = 8'd243; b = 8'd122;  #10 
a = 8'd243; b = 8'd123;  #10 
a = 8'd243; b = 8'd124;  #10 
a = 8'd243; b = 8'd125;  #10 
a = 8'd243; b = 8'd126;  #10 
a = 8'd243; b = 8'd127;  #10 
a = 8'd243; b = 8'd128;  #10 
a = 8'd243; b = 8'd129;  #10 
a = 8'd243; b = 8'd130;  #10 
a = 8'd243; b = 8'd131;  #10 
a = 8'd243; b = 8'd132;  #10 
a = 8'd243; b = 8'd133;  #10 
a = 8'd243; b = 8'd134;  #10 
a = 8'd243; b = 8'd135;  #10 
a = 8'd243; b = 8'd136;  #10 
a = 8'd243; b = 8'd137;  #10 
a = 8'd243; b = 8'd138;  #10 
a = 8'd243; b = 8'd139;  #10 
a = 8'd243; b = 8'd140;  #10 
a = 8'd243; b = 8'd141;  #10 
a = 8'd243; b = 8'd142;  #10 
a = 8'd243; b = 8'd143;  #10 
a = 8'd243; b = 8'd144;  #10 
a = 8'd243; b = 8'd145;  #10 
a = 8'd243; b = 8'd146;  #10 
a = 8'd243; b = 8'd147;  #10 
a = 8'd243; b = 8'd148;  #10 
a = 8'd243; b = 8'd149;  #10 
a = 8'd243; b = 8'd150;  #10 
a = 8'd243; b = 8'd151;  #10 
a = 8'd243; b = 8'd152;  #10 
a = 8'd243; b = 8'd153;  #10 
a = 8'd243; b = 8'd154;  #10 
a = 8'd243; b = 8'd155;  #10 
a = 8'd243; b = 8'd156;  #10 
a = 8'd243; b = 8'd157;  #10 
a = 8'd243; b = 8'd158;  #10 
a = 8'd243; b = 8'd159;  #10 
a = 8'd243; b = 8'd160;  #10 
a = 8'd243; b = 8'd161;  #10 
a = 8'd243; b = 8'd162;  #10 
a = 8'd243; b = 8'd163;  #10 
a = 8'd243; b = 8'd164;  #10 
a = 8'd243; b = 8'd165;  #10 
a = 8'd243; b = 8'd166;  #10 
a = 8'd243; b = 8'd167;  #10 
a = 8'd243; b = 8'd168;  #10 
a = 8'd243; b = 8'd169;  #10 
a = 8'd243; b = 8'd170;  #10 
a = 8'd243; b = 8'd171;  #10 
a = 8'd243; b = 8'd172;  #10 
a = 8'd243; b = 8'd173;  #10 
a = 8'd243; b = 8'd174;  #10 
a = 8'd243; b = 8'd175;  #10 
a = 8'd243; b = 8'd176;  #10 
a = 8'd243; b = 8'd177;  #10 
a = 8'd243; b = 8'd178;  #10 
a = 8'd243; b = 8'd179;  #10 
a = 8'd243; b = 8'd180;  #10 
a = 8'd243; b = 8'd181;  #10 
a = 8'd243; b = 8'd182;  #10 
a = 8'd243; b = 8'd183;  #10 
a = 8'd243; b = 8'd184;  #10 
a = 8'd243; b = 8'd185;  #10 
a = 8'd243; b = 8'd186;  #10 
a = 8'd243; b = 8'd187;  #10 
a = 8'd243; b = 8'd188;  #10 
a = 8'd243; b = 8'd189;  #10 
a = 8'd243; b = 8'd190;  #10 
a = 8'd243; b = 8'd191;  #10 
a = 8'd243; b = 8'd192;  #10 
a = 8'd243; b = 8'd193;  #10 
a = 8'd243; b = 8'd194;  #10 
a = 8'd243; b = 8'd195;  #10 
a = 8'd243; b = 8'd196;  #10 
a = 8'd243; b = 8'd197;  #10 
a = 8'd243; b = 8'd198;  #10 
a = 8'd243; b = 8'd199;  #10 
a = 8'd243; b = 8'd200;  #10 
a = 8'd243; b = 8'd201;  #10 
a = 8'd243; b = 8'd202;  #10 
a = 8'd243; b = 8'd203;  #10 
a = 8'd243; b = 8'd204;  #10 
a = 8'd243; b = 8'd205;  #10 
a = 8'd243; b = 8'd206;  #10 
a = 8'd243; b = 8'd207;  #10 
a = 8'd243; b = 8'd208;  #10 
a = 8'd243; b = 8'd209;  #10 
a = 8'd243; b = 8'd210;  #10 
a = 8'd243; b = 8'd211;  #10 
a = 8'd243; b = 8'd212;  #10 
a = 8'd243; b = 8'd213;  #10 
a = 8'd243; b = 8'd214;  #10 
a = 8'd243; b = 8'd215;  #10 
a = 8'd243; b = 8'd216;  #10 
a = 8'd243; b = 8'd217;  #10 
a = 8'd243; b = 8'd218;  #10 
a = 8'd243; b = 8'd219;  #10 
a = 8'd243; b = 8'd220;  #10 
a = 8'd243; b = 8'd221;  #10 
a = 8'd243; b = 8'd222;  #10 
a = 8'd243; b = 8'd223;  #10 
a = 8'd243; b = 8'd224;  #10 
a = 8'd243; b = 8'd225;  #10 
a = 8'd243; b = 8'd226;  #10 
a = 8'd243; b = 8'd227;  #10 
a = 8'd243; b = 8'd228;  #10 
a = 8'd243; b = 8'd229;  #10 
a = 8'd243; b = 8'd230;  #10 
a = 8'd243; b = 8'd231;  #10 
a = 8'd243; b = 8'd232;  #10 
a = 8'd243; b = 8'd233;  #10 
a = 8'd243; b = 8'd234;  #10 
a = 8'd243; b = 8'd235;  #10 
a = 8'd243; b = 8'd236;  #10 
a = 8'd243; b = 8'd237;  #10 
a = 8'd243; b = 8'd238;  #10 
a = 8'd243; b = 8'd239;  #10 
a = 8'd243; b = 8'd240;  #10 
a = 8'd243; b = 8'd241;  #10 
a = 8'd243; b = 8'd242;  #10 
a = 8'd243; b = 8'd243;  #10 
a = 8'd243; b = 8'd244;  #10 
a = 8'd243; b = 8'd245;  #10 
a = 8'd243; b = 8'd246;  #10 
a = 8'd243; b = 8'd247;  #10 
a = 8'd243; b = 8'd248;  #10 
a = 8'd243; b = 8'd249;  #10 
a = 8'd243; b = 8'd250;  #10 
a = 8'd243; b = 8'd251;  #10 
a = 8'd243; b = 8'd252;  #10 
a = 8'd243; b = 8'd253;  #10 
a = 8'd243; b = 8'd254;  #10 
a = 8'd243; b = 8'd255;  #10 
a = 8'd244; b = 8'd0;  #10 
a = 8'd244; b = 8'd1;  #10 
a = 8'd244; b = 8'd2;  #10 
a = 8'd244; b = 8'd3;  #10 
a = 8'd244; b = 8'd4;  #10 
a = 8'd244; b = 8'd5;  #10 
a = 8'd244; b = 8'd6;  #10 
a = 8'd244; b = 8'd7;  #10 
a = 8'd244; b = 8'd8;  #10 
a = 8'd244; b = 8'd9;  #10 
a = 8'd244; b = 8'd10;  #10 
a = 8'd244; b = 8'd11;  #10 
a = 8'd244; b = 8'd12;  #10 
a = 8'd244; b = 8'd13;  #10 
a = 8'd244; b = 8'd14;  #10 
a = 8'd244; b = 8'd15;  #10 
a = 8'd244; b = 8'd16;  #10 
a = 8'd244; b = 8'd17;  #10 
a = 8'd244; b = 8'd18;  #10 
a = 8'd244; b = 8'd19;  #10 
a = 8'd244; b = 8'd20;  #10 
a = 8'd244; b = 8'd21;  #10 
a = 8'd244; b = 8'd22;  #10 
a = 8'd244; b = 8'd23;  #10 
a = 8'd244; b = 8'd24;  #10 
a = 8'd244; b = 8'd25;  #10 
a = 8'd244; b = 8'd26;  #10 
a = 8'd244; b = 8'd27;  #10 
a = 8'd244; b = 8'd28;  #10 
a = 8'd244; b = 8'd29;  #10 
a = 8'd244; b = 8'd30;  #10 
a = 8'd244; b = 8'd31;  #10 
a = 8'd244; b = 8'd32;  #10 
a = 8'd244; b = 8'd33;  #10 
a = 8'd244; b = 8'd34;  #10 
a = 8'd244; b = 8'd35;  #10 
a = 8'd244; b = 8'd36;  #10 
a = 8'd244; b = 8'd37;  #10 
a = 8'd244; b = 8'd38;  #10 
a = 8'd244; b = 8'd39;  #10 
a = 8'd244; b = 8'd40;  #10 
a = 8'd244; b = 8'd41;  #10 
a = 8'd244; b = 8'd42;  #10 
a = 8'd244; b = 8'd43;  #10 
a = 8'd244; b = 8'd44;  #10 
a = 8'd244; b = 8'd45;  #10 
a = 8'd244; b = 8'd46;  #10 
a = 8'd244; b = 8'd47;  #10 
a = 8'd244; b = 8'd48;  #10 
a = 8'd244; b = 8'd49;  #10 
a = 8'd244; b = 8'd50;  #10 
a = 8'd244; b = 8'd51;  #10 
a = 8'd244; b = 8'd52;  #10 
a = 8'd244; b = 8'd53;  #10 
a = 8'd244; b = 8'd54;  #10 
a = 8'd244; b = 8'd55;  #10 
a = 8'd244; b = 8'd56;  #10 
a = 8'd244; b = 8'd57;  #10 
a = 8'd244; b = 8'd58;  #10 
a = 8'd244; b = 8'd59;  #10 
a = 8'd244; b = 8'd60;  #10 
a = 8'd244; b = 8'd61;  #10 
a = 8'd244; b = 8'd62;  #10 
a = 8'd244; b = 8'd63;  #10 
a = 8'd244; b = 8'd64;  #10 
a = 8'd244; b = 8'd65;  #10 
a = 8'd244; b = 8'd66;  #10 
a = 8'd244; b = 8'd67;  #10 
a = 8'd244; b = 8'd68;  #10 
a = 8'd244; b = 8'd69;  #10 
a = 8'd244; b = 8'd70;  #10 
a = 8'd244; b = 8'd71;  #10 
a = 8'd244; b = 8'd72;  #10 
a = 8'd244; b = 8'd73;  #10 
a = 8'd244; b = 8'd74;  #10 
a = 8'd244; b = 8'd75;  #10 
a = 8'd244; b = 8'd76;  #10 
a = 8'd244; b = 8'd77;  #10 
a = 8'd244; b = 8'd78;  #10 
a = 8'd244; b = 8'd79;  #10 
a = 8'd244; b = 8'd80;  #10 
a = 8'd244; b = 8'd81;  #10 
a = 8'd244; b = 8'd82;  #10 
a = 8'd244; b = 8'd83;  #10 
a = 8'd244; b = 8'd84;  #10 
a = 8'd244; b = 8'd85;  #10 
a = 8'd244; b = 8'd86;  #10 
a = 8'd244; b = 8'd87;  #10 
a = 8'd244; b = 8'd88;  #10 
a = 8'd244; b = 8'd89;  #10 
a = 8'd244; b = 8'd90;  #10 
a = 8'd244; b = 8'd91;  #10 
a = 8'd244; b = 8'd92;  #10 
a = 8'd244; b = 8'd93;  #10 
a = 8'd244; b = 8'd94;  #10 
a = 8'd244; b = 8'd95;  #10 
a = 8'd244; b = 8'd96;  #10 
a = 8'd244; b = 8'd97;  #10 
a = 8'd244; b = 8'd98;  #10 
a = 8'd244; b = 8'd99;  #10 
a = 8'd244; b = 8'd100;  #10 
a = 8'd244; b = 8'd101;  #10 
a = 8'd244; b = 8'd102;  #10 
a = 8'd244; b = 8'd103;  #10 
a = 8'd244; b = 8'd104;  #10 
a = 8'd244; b = 8'd105;  #10 
a = 8'd244; b = 8'd106;  #10 
a = 8'd244; b = 8'd107;  #10 
a = 8'd244; b = 8'd108;  #10 
a = 8'd244; b = 8'd109;  #10 
a = 8'd244; b = 8'd110;  #10 
a = 8'd244; b = 8'd111;  #10 
a = 8'd244; b = 8'd112;  #10 
a = 8'd244; b = 8'd113;  #10 
a = 8'd244; b = 8'd114;  #10 
a = 8'd244; b = 8'd115;  #10 
a = 8'd244; b = 8'd116;  #10 
a = 8'd244; b = 8'd117;  #10 
a = 8'd244; b = 8'd118;  #10 
a = 8'd244; b = 8'd119;  #10 
a = 8'd244; b = 8'd120;  #10 
a = 8'd244; b = 8'd121;  #10 
a = 8'd244; b = 8'd122;  #10 
a = 8'd244; b = 8'd123;  #10 
a = 8'd244; b = 8'd124;  #10 
a = 8'd244; b = 8'd125;  #10 
a = 8'd244; b = 8'd126;  #10 
a = 8'd244; b = 8'd127;  #10 
a = 8'd244; b = 8'd128;  #10 
a = 8'd244; b = 8'd129;  #10 
a = 8'd244; b = 8'd130;  #10 
a = 8'd244; b = 8'd131;  #10 
a = 8'd244; b = 8'd132;  #10 
a = 8'd244; b = 8'd133;  #10 
a = 8'd244; b = 8'd134;  #10 
a = 8'd244; b = 8'd135;  #10 
a = 8'd244; b = 8'd136;  #10 
a = 8'd244; b = 8'd137;  #10 
a = 8'd244; b = 8'd138;  #10 
a = 8'd244; b = 8'd139;  #10 
a = 8'd244; b = 8'd140;  #10 
a = 8'd244; b = 8'd141;  #10 
a = 8'd244; b = 8'd142;  #10 
a = 8'd244; b = 8'd143;  #10 
a = 8'd244; b = 8'd144;  #10 
a = 8'd244; b = 8'd145;  #10 
a = 8'd244; b = 8'd146;  #10 
a = 8'd244; b = 8'd147;  #10 
a = 8'd244; b = 8'd148;  #10 
a = 8'd244; b = 8'd149;  #10 
a = 8'd244; b = 8'd150;  #10 
a = 8'd244; b = 8'd151;  #10 
a = 8'd244; b = 8'd152;  #10 
a = 8'd244; b = 8'd153;  #10 
a = 8'd244; b = 8'd154;  #10 
a = 8'd244; b = 8'd155;  #10 
a = 8'd244; b = 8'd156;  #10 
a = 8'd244; b = 8'd157;  #10 
a = 8'd244; b = 8'd158;  #10 
a = 8'd244; b = 8'd159;  #10 
a = 8'd244; b = 8'd160;  #10 
a = 8'd244; b = 8'd161;  #10 
a = 8'd244; b = 8'd162;  #10 
a = 8'd244; b = 8'd163;  #10 
a = 8'd244; b = 8'd164;  #10 
a = 8'd244; b = 8'd165;  #10 
a = 8'd244; b = 8'd166;  #10 
a = 8'd244; b = 8'd167;  #10 
a = 8'd244; b = 8'd168;  #10 
a = 8'd244; b = 8'd169;  #10 
a = 8'd244; b = 8'd170;  #10 
a = 8'd244; b = 8'd171;  #10 
a = 8'd244; b = 8'd172;  #10 
a = 8'd244; b = 8'd173;  #10 
a = 8'd244; b = 8'd174;  #10 
a = 8'd244; b = 8'd175;  #10 
a = 8'd244; b = 8'd176;  #10 
a = 8'd244; b = 8'd177;  #10 
a = 8'd244; b = 8'd178;  #10 
a = 8'd244; b = 8'd179;  #10 
a = 8'd244; b = 8'd180;  #10 
a = 8'd244; b = 8'd181;  #10 
a = 8'd244; b = 8'd182;  #10 
a = 8'd244; b = 8'd183;  #10 
a = 8'd244; b = 8'd184;  #10 
a = 8'd244; b = 8'd185;  #10 
a = 8'd244; b = 8'd186;  #10 
a = 8'd244; b = 8'd187;  #10 
a = 8'd244; b = 8'd188;  #10 
a = 8'd244; b = 8'd189;  #10 
a = 8'd244; b = 8'd190;  #10 
a = 8'd244; b = 8'd191;  #10 
a = 8'd244; b = 8'd192;  #10 
a = 8'd244; b = 8'd193;  #10 
a = 8'd244; b = 8'd194;  #10 
a = 8'd244; b = 8'd195;  #10 
a = 8'd244; b = 8'd196;  #10 
a = 8'd244; b = 8'd197;  #10 
a = 8'd244; b = 8'd198;  #10 
a = 8'd244; b = 8'd199;  #10 
a = 8'd244; b = 8'd200;  #10 
a = 8'd244; b = 8'd201;  #10 
a = 8'd244; b = 8'd202;  #10 
a = 8'd244; b = 8'd203;  #10 
a = 8'd244; b = 8'd204;  #10 
a = 8'd244; b = 8'd205;  #10 
a = 8'd244; b = 8'd206;  #10 
a = 8'd244; b = 8'd207;  #10 
a = 8'd244; b = 8'd208;  #10 
a = 8'd244; b = 8'd209;  #10 
a = 8'd244; b = 8'd210;  #10 
a = 8'd244; b = 8'd211;  #10 
a = 8'd244; b = 8'd212;  #10 
a = 8'd244; b = 8'd213;  #10 
a = 8'd244; b = 8'd214;  #10 
a = 8'd244; b = 8'd215;  #10 
a = 8'd244; b = 8'd216;  #10 
a = 8'd244; b = 8'd217;  #10 
a = 8'd244; b = 8'd218;  #10 
a = 8'd244; b = 8'd219;  #10 
a = 8'd244; b = 8'd220;  #10 
a = 8'd244; b = 8'd221;  #10 
a = 8'd244; b = 8'd222;  #10 
a = 8'd244; b = 8'd223;  #10 
a = 8'd244; b = 8'd224;  #10 
a = 8'd244; b = 8'd225;  #10 
a = 8'd244; b = 8'd226;  #10 
a = 8'd244; b = 8'd227;  #10 
a = 8'd244; b = 8'd228;  #10 
a = 8'd244; b = 8'd229;  #10 
a = 8'd244; b = 8'd230;  #10 
a = 8'd244; b = 8'd231;  #10 
a = 8'd244; b = 8'd232;  #10 
a = 8'd244; b = 8'd233;  #10 
a = 8'd244; b = 8'd234;  #10 
a = 8'd244; b = 8'd235;  #10 
a = 8'd244; b = 8'd236;  #10 
a = 8'd244; b = 8'd237;  #10 
a = 8'd244; b = 8'd238;  #10 
a = 8'd244; b = 8'd239;  #10 
a = 8'd244; b = 8'd240;  #10 
a = 8'd244; b = 8'd241;  #10 
a = 8'd244; b = 8'd242;  #10 
a = 8'd244; b = 8'd243;  #10 
a = 8'd244; b = 8'd244;  #10 
a = 8'd244; b = 8'd245;  #10 
a = 8'd244; b = 8'd246;  #10 
a = 8'd244; b = 8'd247;  #10 
a = 8'd244; b = 8'd248;  #10 
a = 8'd244; b = 8'd249;  #10 
a = 8'd244; b = 8'd250;  #10 
a = 8'd244; b = 8'd251;  #10 
a = 8'd244; b = 8'd252;  #10 
a = 8'd244; b = 8'd253;  #10 
a = 8'd244; b = 8'd254;  #10 
a = 8'd244; b = 8'd255;  #10 
a = 8'd245; b = 8'd0;  #10 
a = 8'd245; b = 8'd1;  #10 
a = 8'd245; b = 8'd2;  #10 
a = 8'd245; b = 8'd3;  #10 
a = 8'd245; b = 8'd4;  #10 
a = 8'd245; b = 8'd5;  #10 
a = 8'd245; b = 8'd6;  #10 
a = 8'd245; b = 8'd7;  #10 
a = 8'd245; b = 8'd8;  #10 
a = 8'd245; b = 8'd9;  #10 
a = 8'd245; b = 8'd10;  #10 
a = 8'd245; b = 8'd11;  #10 
a = 8'd245; b = 8'd12;  #10 
a = 8'd245; b = 8'd13;  #10 
a = 8'd245; b = 8'd14;  #10 
a = 8'd245; b = 8'd15;  #10 
a = 8'd245; b = 8'd16;  #10 
a = 8'd245; b = 8'd17;  #10 
a = 8'd245; b = 8'd18;  #10 
a = 8'd245; b = 8'd19;  #10 
a = 8'd245; b = 8'd20;  #10 
a = 8'd245; b = 8'd21;  #10 
a = 8'd245; b = 8'd22;  #10 
a = 8'd245; b = 8'd23;  #10 
a = 8'd245; b = 8'd24;  #10 
a = 8'd245; b = 8'd25;  #10 
a = 8'd245; b = 8'd26;  #10 
a = 8'd245; b = 8'd27;  #10 
a = 8'd245; b = 8'd28;  #10 
a = 8'd245; b = 8'd29;  #10 
a = 8'd245; b = 8'd30;  #10 
a = 8'd245; b = 8'd31;  #10 
a = 8'd245; b = 8'd32;  #10 
a = 8'd245; b = 8'd33;  #10 
a = 8'd245; b = 8'd34;  #10 
a = 8'd245; b = 8'd35;  #10 
a = 8'd245; b = 8'd36;  #10 
a = 8'd245; b = 8'd37;  #10 
a = 8'd245; b = 8'd38;  #10 
a = 8'd245; b = 8'd39;  #10 
a = 8'd245; b = 8'd40;  #10 
a = 8'd245; b = 8'd41;  #10 
a = 8'd245; b = 8'd42;  #10 
a = 8'd245; b = 8'd43;  #10 
a = 8'd245; b = 8'd44;  #10 
a = 8'd245; b = 8'd45;  #10 
a = 8'd245; b = 8'd46;  #10 
a = 8'd245; b = 8'd47;  #10 
a = 8'd245; b = 8'd48;  #10 
a = 8'd245; b = 8'd49;  #10 
a = 8'd245; b = 8'd50;  #10 
a = 8'd245; b = 8'd51;  #10 
a = 8'd245; b = 8'd52;  #10 
a = 8'd245; b = 8'd53;  #10 
a = 8'd245; b = 8'd54;  #10 
a = 8'd245; b = 8'd55;  #10 
a = 8'd245; b = 8'd56;  #10 
a = 8'd245; b = 8'd57;  #10 
a = 8'd245; b = 8'd58;  #10 
a = 8'd245; b = 8'd59;  #10 
a = 8'd245; b = 8'd60;  #10 
a = 8'd245; b = 8'd61;  #10 
a = 8'd245; b = 8'd62;  #10 
a = 8'd245; b = 8'd63;  #10 
a = 8'd245; b = 8'd64;  #10 
a = 8'd245; b = 8'd65;  #10 
a = 8'd245; b = 8'd66;  #10 
a = 8'd245; b = 8'd67;  #10 
a = 8'd245; b = 8'd68;  #10 
a = 8'd245; b = 8'd69;  #10 
a = 8'd245; b = 8'd70;  #10 
a = 8'd245; b = 8'd71;  #10 
a = 8'd245; b = 8'd72;  #10 
a = 8'd245; b = 8'd73;  #10 
a = 8'd245; b = 8'd74;  #10 
a = 8'd245; b = 8'd75;  #10 
a = 8'd245; b = 8'd76;  #10 
a = 8'd245; b = 8'd77;  #10 
a = 8'd245; b = 8'd78;  #10 
a = 8'd245; b = 8'd79;  #10 
a = 8'd245; b = 8'd80;  #10 
a = 8'd245; b = 8'd81;  #10 
a = 8'd245; b = 8'd82;  #10 
a = 8'd245; b = 8'd83;  #10 
a = 8'd245; b = 8'd84;  #10 
a = 8'd245; b = 8'd85;  #10 
a = 8'd245; b = 8'd86;  #10 
a = 8'd245; b = 8'd87;  #10 
a = 8'd245; b = 8'd88;  #10 
a = 8'd245; b = 8'd89;  #10 
a = 8'd245; b = 8'd90;  #10 
a = 8'd245; b = 8'd91;  #10 
a = 8'd245; b = 8'd92;  #10 
a = 8'd245; b = 8'd93;  #10 
a = 8'd245; b = 8'd94;  #10 
a = 8'd245; b = 8'd95;  #10 
a = 8'd245; b = 8'd96;  #10 
a = 8'd245; b = 8'd97;  #10 
a = 8'd245; b = 8'd98;  #10 
a = 8'd245; b = 8'd99;  #10 
a = 8'd245; b = 8'd100;  #10 
a = 8'd245; b = 8'd101;  #10 
a = 8'd245; b = 8'd102;  #10 
a = 8'd245; b = 8'd103;  #10 
a = 8'd245; b = 8'd104;  #10 
a = 8'd245; b = 8'd105;  #10 
a = 8'd245; b = 8'd106;  #10 
a = 8'd245; b = 8'd107;  #10 
a = 8'd245; b = 8'd108;  #10 
a = 8'd245; b = 8'd109;  #10 
a = 8'd245; b = 8'd110;  #10 
a = 8'd245; b = 8'd111;  #10 
a = 8'd245; b = 8'd112;  #10 
a = 8'd245; b = 8'd113;  #10 
a = 8'd245; b = 8'd114;  #10 
a = 8'd245; b = 8'd115;  #10 
a = 8'd245; b = 8'd116;  #10 
a = 8'd245; b = 8'd117;  #10 
a = 8'd245; b = 8'd118;  #10 
a = 8'd245; b = 8'd119;  #10 
a = 8'd245; b = 8'd120;  #10 
a = 8'd245; b = 8'd121;  #10 
a = 8'd245; b = 8'd122;  #10 
a = 8'd245; b = 8'd123;  #10 
a = 8'd245; b = 8'd124;  #10 
a = 8'd245; b = 8'd125;  #10 
a = 8'd245; b = 8'd126;  #10 
a = 8'd245; b = 8'd127;  #10 
a = 8'd245; b = 8'd128;  #10 
a = 8'd245; b = 8'd129;  #10 
a = 8'd245; b = 8'd130;  #10 
a = 8'd245; b = 8'd131;  #10 
a = 8'd245; b = 8'd132;  #10 
a = 8'd245; b = 8'd133;  #10 
a = 8'd245; b = 8'd134;  #10 
a = 8'd245; b = 8'd135;  #10 
a = 8'd245; b = 8'd136;  #10 
a = 8'd245; b = 8'd137;  #10 
a = 8'd245; b = 8'd138;  #10 
a = 8'd245; b = 8'd139;  #10 
a = 8'd245; b = 8'd140;  #10 
a = 8'd245; b = 8'd141;  #10 
a = 8'd245; b = 8'd142;  #10 
a = 8'd245; b = 8'd143;  #10 
a = 8'd245; b = 8'd144;  #10 
a = 8'd245; b = 8'd145;  #10 
a = 8'd245; b = 8'd146;  #10 
a = 8'd245; b = 8'd147;  #10 
a = 8'd245; b = 8'd148;  #10 
a = 8'd245; b = 8'd149;  #10 
a = 8'd245; b = 8'd150;  #10 
a = 8'd245; b = 8'd151;  #10 
a = 8'd245; b = 8'd152;  #10 
a = 8'd245; b = 8'd153;  #10 
a = 8'd245; b = 8'd154;  #10 
a = 8'd245; b = 8'd155;  #10 
a = 8'd245; b = 8'd156;  #10 
a = 8'd245; b = 8'd157;  #10 
a = 8'd245; b = 8'd158;  #10 
a = 8'd245; b = 8'd159;  #10 
a = 8'd245; b = 8'd160;  #10 
a = 8'd245; b = 8'd161;  #10 
a = 8'd245; b = 8'd162;  #10 
a = 8'd245; b = 8'd163;  #10 
a = 8'd245; b = 8'd164;  #10 
a = 8'd245; b = 8'd165;  #10 
a = 8'd245; b = 8'd166;  #10 
a = 8'd245; b = 8'd167;  #10 
a = 8'd245; b = 8'd168;  #10 
a = 8'd245; b = 8'd169;  #10 
a = 8'd245; b = 8'd170;  #10 
a = 8'd245; b = 8'd171;  #10 
a = 8'd245; b = 8'd172;  #10 
a = 8'd245; b = 8'd173;  #10 
a = 8'd245; b = 8'd174;  #10 
a = 8'd245; b = 8'd175;  #10 
a = 8'd245; b = 8'd176;  #10 
a = 8'd245; b = 8'd177;  #10 
a = 8'd245; b = 8'd178;  #10 
a = 8'd245; b = 8'd179;  #10 
a = 8'd245; b = 8'd180;  #10 
a = 8'd245; b = 8'd181;  #10 
a = 8'd245; b = 8'd182;  #10 
a = 8'd245; b = 8'd183;  #10 
a = 8'd245; b = 8'd184;  #10 
a = 8'd245; b = 8'd185;  #10 
a = 8'd245; b = 8'd186;  #10 
a = 8'd245; b = 8'd187;  #10 
a = 8'd245; b = 8'd188;  #10 
a = 8'd245; b = 8'd189;  #10 
a = 8'd245; b = 8'd190;  #10 
a = 8'd245; b = 8'd191;  #10 
a = 8'd245; b = 8'd192;  #10 
a = 8'd245; b = 8'd193;  #10 
a = 8'd245; b = 8'd194;  #10 
a = 8'd245; b = 8'd195;  #10 
a = 8'd245; b = 8'd196;  #10 
a = 8'd245; b = 8'd197;  #10 
a = 8'd245; b = 8'd198;  #10 
a = 8'd245; b = 8'd199;  #10 
a = 8'd245; b = 8'd200;  #10 
a = 8'd245; b = 8'd201;  #10 
a = 8'd245; b = 8'd202;  #10 
a = 8'd245; b = 8'd203;  #10 
a = 8'd245; b = 8'd204;  #10 
a = 8'd245; b = 8'd205;  #10 
a = 8'd245; b = 8'd206;  #10 
a = 8'd245; b = 8'd207;  #10 
a = 8'd245; b = 8'd208;  #10 
a = 8'd245; b = 8'd209;  #10 
a = 8'd245; b = 8'd210;  #10 
a = 8'd245; b = 8'd211;  #10 
a = 8'd245; b = 8'd212;  #10 
a = 8'd245; b = 8'd213;  #10 
a = 8'd245; b = 8'd214;  #10 
a = 8'd245; b = 8'd215;  #10 
a = 8'd245; b = 8'd216;  #10 
a = 8'd245; b = 8'd217;  #10 
a = 8'd245; b = 8'd218;  #10 
a = 8'd245; b = 8'd219;  #10 
a = 8'd245; b = 8'd220;  #10 
a = 8'd245; b = 8'd221;  #10 
a = 8'd245; b = 8'd222;  #10 
a = 8'd245; b = 8'd223;  #10 
a = 8'd245; b = 8'd224;  #10 
a = 8'd245; b = 8'd225;  #10 
a = 8'd245; b = 8'd226;  #10 
a = 8'd245; b = 8'd227;  #10 
a = 8'd245; b = 8'd228;  #10 
a = 8'd245; b = 8'd229;  #10 
a = 8'd245; b = 8'd230;  #10 
a = 8'd245; b = 8'd231;  #10 
a = 8'd245; b = 8'd232;  #10 
a = 8'd245; b = 8'd233;  #10 
a = 8'd245; b = 8'd234;  #10 
a = 8'd245; b = 8'd235;  #10 
a = 8'd245; b = 8'd236;  #10 
a = 8'd245; b = 8'd237;  #10 
a = 8'd245; b = 8'd238;  #10 
a = 8'd245; b = 8'd239;  #10 
a = 8'd245; b = 8'd240;  #10 
a = 8'd245; b = 8'd241;  #10 
a = 8'd245; b = 8'd242;  #10 
a = 8'd245; b = 8'd243;  #10 
a = 8'd245; b = 8'd244;  #10 
a = 8'd245; b = 8'd245;  #10 
a = 8'd245; b = 8'd246;  #10 
a = 8'd245; b = 8'd247;  #10 
a = 8'd245; b = 8'd248;  #10 
a = 8'd245; b = 8'd249;  #10 
a = 8'd245; b = 8'd250;  #10 
a = 8'd245; b = 8'd251;  #10 
a = 8'd245; b = 8'd252;  #10 
a = 8'd245; b = 8'd253;  #10 
a = 8'd245; b = 8'd254;  #10 
a = 8'd245; b = 8'd255;  #10 
a = 8'd246; b = 8'd0;  #10 
a = 8'd246; b = 8'd1;  #10 
a = 8'd246; b = 8'd2;  #10 
a = 8'd246; b = 8'd3;  #10 
a = 8'd246; b = 8'd4;  #10 
a = 8'd246; b = 8'd5;  #10 
a = 8'd246; b = 8'd6;  #10 
a = 8'd246; b = 8'd7;  #10 
a = 8'd246; b = 8'd8;  #10 
a = 8'd246; b = 8'd9;  #10 
a = 8'd246; b = 8'd10;  #10 
a = 8'd246; b = 8'd11;  #10 
a = 8'd246; b = 8'd12;  #10 
a = 8'd246; b = 8'd13;  #10 
a = 8'd246; b = 8'd14;  #10 
a = 8'd246; b = 8'd15;  #10 
a = 8'd246; b = 8'd16;  #10 
a = 8'd246; b = 8'd17;  #10 
a = 8'd246; b = 8'd18;  #10 
a = 8'd246; b = 8'd19;  #10 
a = 8'd246; b = 8'd20;  #10 
a = 8'd246; b = 8'd21;  #10 
a = 8'd246; b = 8'd22;  #10 
a = 8'd246; b = 8'd23;  #10 
a = 8'd246; b = 8'd24;  #10 
a = 8'd246; b = 8'd25;  #10 
a = 8'd246; b = 8'd26;  #10 
a = 8'd246; b = 8'd27;  #10 
a = 8'd246; b = 8'd28;  #10 
a = 8'd246; b = 8'd29;  #10 
a = 8'd246; b = 8'd30;  #10 
a = 8'd246; b = 8'd31;  #10 
a = 8'd246; b = 8'd32;  #10 
a = 8'd246; b = 8'd33;  #10 
a = 8'd246; b = 8'd34;  #10 
a = 8'd246; b = 8'd35;  #10 
a = 8'd246; b = 8'd36;  #10 
a = 8'd246; b = 8'd37;  #10 
a = 8'd246; b = 8'd38;  #10 
a = 8'd246; b = 8'd39;  #10 
a = 8'd246; b = 8'd40;  #10 
a = 8'd246; b = 8'd41;  #10 
a = 8'd246; b = 8'd42;  #10 
a = 8'd246; b = 8'd43;  #10 
a = 8'd246; b = 8'd44;  #10 
a = 8'd246; b = 8'd45;  #10 
a = 8'd246; b = 8'd46;  #10 
a = 8'd246; b = 8'd47;  #10 
a = 8'd246; b = 8'd48;  #10 
a = 8'd246; b = 8'd49;  #10 
a = 8'd246; b = 8'd50;  #10 
a = 8'd246; b = 8'd51;  #10 
a = 8'd246; b = 8'd52;  #10 
a = 8'd246; b = 8'd53;  #10 
a = 8'd246; b = 8'd54;  #10 
a = 8'd246; b = 8'd55;  #10 
a = 8'd246; b = 8'd56;  #10 
a = 8'd246; b = 8'd57;  #10 
a = 8'd246; b = 8'd58;  #10 
a = 8'd246; b = 8'd59;  #10 
a = 8'd246; b = 8'd60;  #10 
a = 8'd246; b = 8'd61;  #10 
a = 8'd246; b = 8'd62;  #10 
a = 8'd246; b = 8'd63;  #10 
a = 8'd246; b = 8'd64;  #10 
a = 8'd246; b = 8'd65;  #10 
a = 8'd246; b = 8'd66;  #10 
a = 8'd246; b = 8'd67;  #10 
a = 8'd246; b = 8'd68;  #10 
a = 8'd246; b = 8'd69;  #10 
a = 8'd246; b = 8'd70;  #10 
a = 8'd246; b = 8'd71;  #10 
a = 8'd246; b = 8'd72;  #10 
a = 8'd246; b = 8'd73;  #10 
a = 8'd246; b = 8'd74;  #10 
a = 8'd246; b = 8'd75;  #10 
a = 8'd246; b = 8'd76;  #10 
a = 8'd246; b = 8'd77;  #10 
a = 8'd246; b = 8'd78;  #10 
a = 8'd246; b = 8'd79;  #10 
a = 8'd246; b = 8'd80;  #10 
a = 8'd246; b = 8'd81;  #10 
a = 8'd246; b = 8'd82;  #10 
a = 8'd246; b = 8'd83;  #10 
a = 8'd246; b = 8'd84;  #10 
a = 8'd246; b = 8'd85;  #10 
a = 8'd246; b = 8'd86;  #10 
a = 8'd246; b = 8'd87;  #10 
a = 8'd246; b = 8'd88;  #10 
a = 8'd246; b = 8'd89;  #10 
a = 8'd246; b = 8'd90;  #10 
a = 8'd246; b = 8'd91;  #10 
a = 8'd246; b = 8'd92;  #10 
a = 8'd246; b = 8'd93;  #10 
a = 8'd246; b = 8'd94;  #10 
a = 8'd246; b = 8'd95;  #10 
a = 8'd246; b = 8'd96;  #10 
a = 8'd246; b = 8'd97;  #10 
a = 8'd246; b = 8'd98;  #10 
a = 8'd246; b = 8'd99;  #10 
a = 8'd246; b = 8'd100;  #10 
a = 8'd246; b = 8'd101;  #10 
a = 8'd246; b = 8'd102;  #10 
a = 8'd246; b = 8'd103;  #10 
a = 8'd246; b = 8'd104;  #10 
a = 8'd246; b = 8'd105;  #10 
a = 8'd246; b = 8'd106;  #10 
a = 8'd246; b = 8'd107;  #10 
a = 8'd246; b = 8'd108;  #10 
a = 8'd246; b = 8'd109;  #10 
a = 8'd246; b = 8'd110;  #10 
a = 8'd246; b = 8'd111;  #10 
a = 8'd246; b = 8'd112;  #10 
a = 8'd246; b = 8'd113;  #10 
a = 8'd246; b = 8'd114;  #10 
a = 8'd246; b = 8'd115;  #10 
a = 8'd246; b = 8'd116;  #10 
a = 8'd246; b = 8'd117;  #10 
a = 8'd246; b = 8'd118;  #10 
a = 8'd246; b = 8'd119;  #10 
a = 8'd246; b = 8'd120;  #10 
a = 8'd246; b = 8'd121;  #10 
a = 8'd246; b = 8'd122;  #10 
a = 8'd246; b = 8'd123;  #10 
a = 8'd246; b = 8'd124;  #10 
a = 8'd246; b = 8'd125;  #10 
a = 8'd246; b = 8'd126;  #10 
a = 8'd246; b = 8'd127;  #10 
a = 8'd246; b = 8'd128;  #10 
a = 8'd246; b = 8'd129;  #10 
a = 8'd246; b = 8'd130;  #10 
a = 8'd246; b = 8'd131;  #10 
a = 8'd246; b = 8'd132;  #10 
a = 8'd246; b = 8'd133;  #10 
a = 8'd246; b = 8'd134;  #10 
a = 8'd246; b = 8'd135;  #10 
a = 8'd246; b = 8'd136;  #10 
a = 8'd246; b = 8'd137;  #10 
a = 8'd246; b = 8'd138;  #10 
a = 8'd246; b = 8'd139;  #10 
a = 8'd246; b = 8'd140;  #10 
a = 8'd246; b = 8'd141;  #10 
a = 8'd246; b = 8'd142;  #10 
a = 8'd246; b = 8'd143;  #10 
a = 8'd246; b = 8'd144;  #10 
a = 8'd246; b = 8'd145;  #10 
a = 8'd246; b = 8'd146;  #10 
a = 8'd246; b = 8'd147;  #10 
a = 8'd246; b = 8'd148;  #10 
a = 8'd246; b = 8'd149;  #10 
a = 8'd246; b = 8'd150;  #10 
a = 8'd246; b = 8'd151;  #10 
a = 8'd246; b = 8'd152;  #10 
a = 8'd246; b = 8'd153;  #10 
a = 8'd246; b = 8'd154;  #10 
a = 8'd246; b = 8'd155;  #10 
a = 8'd246; b = 8'd156;  #10 
a = 8'd246; b = 8'd157;  #10 
a = 8'd246; b = 8'd158;  #10 
a = 8'd246; b = 8'd159;  #10 
a = 8'd246; b = 8'd160;  #10 
a = 8'd246; b = 8'd161;  #10 
a = 8'd246; b = 8'd162;  #10 
a = 8'd246; b = 8'd163;  #10 
a = 8'd246; b = 8'd164;  #10 
a = 8'd246; b = 8'd165;  #10 
a = 8'd246; b = 8'd166;  #10 
a = 8'd246; b = 8'd167;  #10 
a = 8'd246; b = 8'd168;  #10 
a = 8'd246; b = 8'd169;  #10 
a = 8'd246; b = 8'd170;  #10 
a = 8'd246; b = 8'd171;  #10 
a = 8'd246; b = 8'd172;  #10 
a = 8'd246; b = 8'd173;  #10 
a = 8'd246; b = 8'd174;  #10 
a = 8'd246; b = 8'd175;  #10 
a = 8'd246; b = 8'd176;  #10 
a = 8'd246; b = 8'd177;  #10 
a = 8'd246; b = 8'd178;  #10 
a = 8'd246; b = 8'd179;  #10 
a = 8'd246; b = 8'd180;  #10 
a = 8'd246; b = 8'd181;  #10 
a = 8'd246; b = 8'd182;  #10 
a = 8'd246; b = 8'd183;  #10 
a = 8'd246; b = 8'd184;  #10 
a = 8'd246; b = 8'd185;  #10 
a = 8'd246; b = 8'd186;  #10 
a = 8'd246; b = 8'd187;  #10 
a = 8'd246; b = 8'd188;  #10 
a = 8'd246; b = 8'd189;  #10 
a = 8'd246; b = 8'd190;  #10 
a = 8'd246; b = 8'd191;  #10 
a = 8'd246; b = 8'd192;  #10 
a = 8'd246; b = 8'd193;  #10 
a = 8'd246; b = 8'd194;  #10 
a = 8'd246; b = 8'd195;  #10 
a = 8'd246; b = 8'd196;  #10 
a = 8'd246; b = 8'd197;  #10 
a = 8'd246; b = 8'd198;  #10 
a = 8'd246; b = 8'd199;  #10 
a = 8'd246; b = 8'd200;  #10 
a = 8'd246; b = 8'd201;  #10 
a = 8'd246; b = 8'd202;  #10 
a = 8'd246; b = 8'd203;  #10 
a = 8'd246; b = 8'd204;  #10 
a = 8'd246; b = 8'd205;  #10 
a = 8'd246; b = 8'd206;  #10 
a = 8'd246; b = 8'd207;  #10 
a = 8'd246; b = 8'd208;  #10 
a = 8'd246; b = 8'd209;  #10 
a = 8'd246; b = 8'd210;  #10 
a = 8'd246; b = 8'd211;  #10 
a = 8'd246; b = 8'd212;  #10 
a = 8'd246; b = 8'd213;  #10 
a = 8'd246; b = 8'd214;  #10 
a = 8'd246; b = 8'd215;  #10 
a = 8'd246; b = 8'd216;  #10 
a = 8'd246; b = 8'd217;  #10 
a = 8'd246; b = 8'd218;  #10 
a = 8'd246; b = 8'd219;  #10 
a = 8'd246; b = 8'd220;  #10 
a = 8'd246; b = 8'd221;  #10 
a = 8'd246; b = 8'd222;  #10 
a = 8'd246; b = 8'd223;  #10 
a = 8'd246; b = 8'd224;  #10 
a = 8'd246; b = 8'd225;  #10 
a = 8'd246; b = 8'd226;  #10 
a = 8'd246; b = 8'd227;  #10 
a = 8'd246; b = 8'd228;  #10 
a = 8'd246; b = 8'd229;  #10 
a = 8'd246; b = 8'd230;  #10 
a = 8'd246; b = 8'd231;  #10 
a = 8'd246; b = 8'd232;  #10 
a = 8'd246; b = 8'd233;  #10 
a = 8'd246; b = 8'd234;  #10 
a = 8'd246; b = 8'd235;  #10 
a = 8'd246; b = 8'd236;  #10 
a = 8'd246; b = 8'd237;  #10 
a = 8'd246; b = 8'd238;  #10 
a = 8'd246; b = 8'd239;  #10 
a = 8'd246; b = 8'd240;  #10 
a = 8'd246; b = 8'd241;  #10 
a = 8'd246; b = 8'd242;  #10 
a = 8'd246; b = 8'd243;  #10 
a = 8'd246; b = 8'd244;  #10 
a = 8'd246; b = 8'd245;  #10 
a = 8'd246; b = 8'd246;  #10 
a = 8'd246; b = 8'd247;  #10 
a = 8'd246; b = 8'd248;  #10 
a = 8'd246; b = 8'd249;  #10 
a = 8'd246; b = 8'd250;  #10 
a = 8'd246; b = 8'd251;  #10 
a = 8'd246; b = 8'd252;  #10 
a = 8'd246; b = 8'd253;  #10 
a = 8'd246; b = 8'd254;  #10 
a = 8'd246; b = 8'd255;  #10 
a = 8'd247; b = 8'd0;  #10 
a = 8'd247; b = 8'd1;  #10 
a = 8'd247; b = 8'd2;  #10 
a = 8'd247; b = 8'd3;  #10 
a = 8'd247; b = 8'd4;  #10 
a = 8'd247; b = 8'd5;  #10 
a = 8'd247; b = 8'd6;  #10 
a = 8'd247; b = 8'd7;  #10 
a = 8'd247; b = 8'd8;  #10 
a = 8'd247; b = 8'd9;  #10 
a = 8'd247; b = 8'd10;  #10 
a = 8'd247; b = 8'd11;  #10 
a = 8'd247; b = 8'd12;  #10 
a = 8'd247; b = 8'd13;  #10 
a = 8'd247; b = 8'd14;  #10 
a = 8'd247; b = 8'd15;  #10 
a = 8'd247; b = 8'd16;  #10 
a = 8'd247; b = 8'd17;  #10 
a = 8'd247; b = 8'd18;  #10 
a = 8'd247; b = 8'd19;  #10 
a = 8'd247; b = 8'd20;  #10 
a = 8'd247; b = 8'd21;  #10 
a = 8'd247; b = 8'd22;  #10 
a = 8'd247; b = 8'd23;  #10 
a = 8'd247; b = 8'd24;  #10 
a = 8'd247; b = 8'd25;  #10 
a = 8'd247; b = 8'd26;  #10 
a = 8'd247; b = 8'd27;  #10 
a = 8'd247; b = 8'd28;  #10 
a = 8'd247; b = 8'd29;  #10 
a = 8'd247; b = 8'd30;  #10 
a = 8'd247; b = 8'd31;  #10 
a = 8'd247; b = 8'd32;  #10 
a = 8'd247; b = 8'd33;  #10 
a = 8'd247; b = 8'd34;  #10 
a = 8'd247; b = 8'd35;  #10 
a = 8'd247; b = 8'd36;  #10 
a = 8'd247; b = 8'd37;  #10 
a = 8'd247; b = 8'd38;  #10 
a = 8'd247; b = 8'd39;  #10 
a = 8'd247; b = 8'd40;  #10 
a = 8'd247; b = 8'd41;  #10 
a = 8'd247; b = 8'd42;  #10 
a = 8'd247; b = 8'd43;  #10 
a = 8'd247; b = 8'd44;  #10 
a = 8'd247; b = 8'd45;  #10 
a = 8'd247; b = 8'd46;  #10 
a = 8'd247; b = 8'd47;  #10 
a = 8'd247; b = 8'd48;  #10 
a = 8'd247; b = 8'd49;  #10 
a = 8'd247; b = 8'd50;  #10 
a = 8'd247; b = 8'd51;  #10 
a = 8'd247; b = 8'd52;  #10 
a = 8'd247; b = 8'd53;  #10 
a = 8'd247; b = 8'd54;  #10 
a = 8'd247; b = 8'd55;  #10 
a = 8'd247; b = 8'd56;  #10 
a = 8'd247; b = 8'd57;  #10 
a = 8'd247; b = 8'd58;  #10 
a = 8'd247; b = 8'd59;  #10 
a = 8'd247; b = 8'd60;  #10 
a = 8'd247; b = 8'd61;  #10 
a = 8'd247; b = 8'd62;  #10 
a = 8'd247; b = 8'd63;  #10 
a = 8'd247; b = 8'd64;  #10 
a = 8'd247; b = 8'd65;  #10 
a = 8'd247; b = 8'd66;  #10 
a = 8'd247; b = 8'd67;  #10 
a = 8'd247; b = 8'd68;  #10 
a = 8'd247; b = 8'd69;  #10 
a = 8'd247; b = 8'd70;  #10 
a = 8'd247; b = 8'd71;  #10 
a = 8'd247; b = 8'd72;  #10 
a = 8'd247; b = 8'd73;  #10 
a = 8'd247; b = 8'd74;  #10 
a = 8'd247; b = 8'd75;  #10 
a = 8'd247; b = 8'd76;  #10 
a = 8'd247; b = 8'd77;  #10 
a = 8'd247; b = 8'd78;  #10 
a = 8'd247; b = 8'd79;  #10 
a = 8'd247; b = 8'd80;  #10 
a = 8'd247; b = 8'd81;  #10 
a = 8'd247; b = 8'd82;  #10 
a = 8'd247; b = 8'd83;  #10 
a = 8'd247; b = 8'd84;  #10 
a = 8'd247; b = 8'd85;  #10 
a = 8'd247; b = 8'd86;  #10 
a = 8'd247; b = 8'd87;  #10 
a = 8'd247; b = 8'd88;  #10 
a = 8'd247; b = 8'd89;  #10 
a = 8'd247; b = 8'd90;  #10 
a = 8'd247; b = 8'd91;  #10 
a = 8'd247; b = 8'd92;  #10 
a = 8'd247; b = 8'd93;  #10 
a = 8'd247; b = 8'd94;  #10 
a = 8'd247; b = 8'd95;  #10 
a = 8'd247; b = 8'd96;  #10 
a = 8'd247; b = 8'd97;  #10 
a = 8'd247; b = 8'd98;  #10 
a = 8'd247; b = 8'd99;  #10 
a = 8'd247; b = 8'd100;  #10 
a = 8'd247; b = 8'd101;  #10 
a = 8'd247; b = 8'd102;  #10 
a = 8'd247; b = 8'd103;  #10 
a = 8'd247; b = 8'd104;  #10 
a = 8'd247; b = 8'd105;  #10 
a = 8'd247; b = 8'd106;  #10 
a = 8'd247; b = 8'd107;  #10 
a = 8'd247; b = 8'd108;  #10 
a = 8'd247; b = 8'd109;  #10 
a = 8'd247; b = 8'd110;  #10 
a = 8'd247; b = 8'd111;  #10 
a = 8'd247; b = 8'd112;  #10 
a = 8'd247; b = 8'd113;  #10 
a = 8'd247; b = 8'd114;  #10 
a = 8'd247; b = 8'd115;  #10 
a = 8'd247; b = 8'd116;  #10 
a = 8'd247; b = 8'd117;  #10 
a = 8'd247; b = 8'd118;  #10 
a = 8'd247; b = 8'd119;  #10 
a = 8'd247; b = 8'd120;  #10 
a = 8'd247; b = 8'd121;  #10 
a = 8'd247; b = 8'd122;  #10 
a = 8'd247; b = 8'd123;  #10 
a = 8'd247; b = 8'd124;  #10 
a = 8'd247; b = 8'd125;  #10 
a = 8'd247; b = 8'd126;  #10 
a = 8'd247; b = 8'd127;  #10 
a = 8'd247; b = 8'd128;  #10 
a = 8'd247; b = 8'd129;  #10 
a = 8'd247; b = 8'd130;  #10 
a = 8'd247; b = 8'd131;  #10 
a = 8'd247; b = 8'd132;  #10 
a = 8'd247; b = 8'd133;  #10 
a = 8'd247; b = 8'd134;  #10 
a = 8'd247; b = 8'd135;  #10 
a = 8'd247; b = 8'd136;  #10 
a = 8'd247; b = 8'd137;  #10 
a = 8'd247; b = 8'd138;  #10 
a = 8'd247; b = 8'd139;  #10 
a = 8'd247; b = 8'd140;  #10 
a = 8'd247; b = 8'd141;  #10 
a = 8'd247; b = 8'd142;  #10 
a = 8'd247; b = 8'd143;  #10 
a = 8'd247; b = 8'd144;  #10 
a = 8'd247; b = 8'd145;  #10 
a = 8'd247; b = 8'd146;  #10 
a = 8'd247; b = 8'd147;  #10 
a = 8'd247; b = 8'd148;  #10 
a = 8'd247; b = 8'd149;  #10 
a = 8'd247; b = 8'd150;  #10 
a = 8'd247; b = 8'd151;  #10 
a = 8'd247; b = 8'd152;  #10 
a = 8'd247; b = 8'd153;  #10 
a = 8'd247; b = 8'd154;  #10 
a = 8'd247; b = 8'd155;  #10 
a = 8'd247; b = 8'd156;  #10 
a = 8'd247; b = 8'd157;  #10 
a = 8'd247; b = 8'd158;  #10 
a = 8'd247; b = 8'd159;  #10 
a = 8'd247; b = 8'd160;  #10 
a = 8'd247; b = 8'd161;  #10 
a = 8'd247; b = 8'd162;  #10 
a = 8'd247; b = 8'd163;  #10 
a = 8'd247; b = 8'd164;  #10 
a = 8'd247; b = 8'd165;  #10 
a = 8'd247; b = 8'd166;  #10 
a = 8'd247; b = 8'd167;  #10 
a = 8'd247; b = 8'd168;  #10 
a = 8'd247; b = 8'd169;  #10 
a = 8'd247; b = 8'd170;  #10 
a = 8'd247; b = 8'd171;  #10 
a = 8'd247; b = 8'd172;  #10 
a = 8'd247; b = 8'd173;  #10 
a = 8'd247; b = 8'd174;  #10 
a = 8'd247; b = 8'd175;  #10 
a = 8'd247; b = 8'd176;  #10 
a = 8'd247; b = 8'd177;  #10 
a = 8'd247; b = 8'd178;  #10 
a = 8'd247; b = 8'd179;  #10 
a = 8'd247; b = 8'd180;  #10 
a = 8'd247; b = 8'd181;  #10 
a = 8'd247; b = 8'd182;  #10 
a = 8'd247; b = 8'd183;  #10 
a = 8'd247; b = 8'd184;  #10 
a = 8'd247; b = 8'd185;  #10 
a = 8'd247; b = 8'd186;  #10 
a = 8'd247; b = 8'd187;  #10 
a = 8'd247; b = 8'd188;  #10 
a = 8'd247; b = 8'd189;  #10 
a = 8'd247; b = 8'd190;  #10 
a = 8'd247; b = 8'd191;  #10 
a = 8'd247; b = 8'd192;  #10 
a = 8'd247; b = 8'd193;  #10 
a = 8'd247; b = 8'd194;  #10 
a = 8'd247; b = 8'd195;  #10 
a = 8'd247; b = 8'd196;  #10 
a = 8'd247; b = 8'd197;  #10 
a = 8'd247; b = 8'd198;  #10 
a = 8'd247; b = 8'd199;  #10 
a = 8'd247; b = 8'd200;  #10 
a = 8'd247; b = 8'd201;  #10 
a = 8'd247; b = 8'd202;  #10 
a = 8'd247; b = 8'd203;  #10 
a = 8'd247; b = 8'd204;  #10 
a = 8'd247; b = 8'd205;  #10 
a = 8'd247; b = 8'd206;  #10 
a = 8'd247; b = 8'd207;  #10 
a = 8'd247; b = 8'd208;  #10 
a = 8'd247; b = 8'd209;  #10 
a = 8'd247; b = 8'd210;  #10 
a = 8'd247; b = 8'd211;  #10 
a = 8'd247; b = 8'd212;  #10 
a = 8'd247; b = 8'd213;  #10 
a = 8'd247; b = 8'd214;  #10 
a = 8'd247; b = 8'd215;  #10 
a = 8'd247; b = 8'd216;  #10 
a = 8'd247; b = 8'd217;  #10 
a = 8'd247; b = 8'd218;  #10 
a = 8'd247; b = 8'd219;  #10 
a = 8'd247; b = 8'd220;  #10 
a = 8'd247; b = 8'd221;  #10 
a = 8'd247; b = 8'd222;  #10 
a = 8'd247; b = 8'd223;  #10 
a = 8'd247; b = 8'd224;  #10 
a = 8'd247; b = 8'd225;  #10 
a = 8'd247; b = 8'd226;  #10 
a = 8'd247; b = 8'd227;  #10 
a = 8'd247; b = 8'd228;  #10 
a = 8'd247; b = 8'd229;  #10 
a = 8'd247; b = 8'd230;  #10 
a = 8'd247; b = 8'd231;  #10 
a = 8'd247; b = 8'd232;  #10 
a = 8'd247; b = 8'd233;  #10 
a = 8'd247; b = 8'd234;  #10 
a = 8'd247; b = 8'd235;  #10 
a = 8'd247; b = 8'd236;  #10 
a = 8'd247; b = 8'd237;  #10 
a = 8'd247; b = 8'd238;  #10 
a = 8'd247; b = 8'd239;  #10 
a = 8'd247; b = 8'd240;  #10 
a = 8'd247; b = 8'd241;  #10 
a = 8'd247; b = 8'd242;  #10 
a = 8'd247; b = 8'd243;  #10 
a = 8'd247; b = 8'd244;  #10 
a = 8'd247; b = 8'd245;  #10 
a = 8'd247; b = 8'd246;  #10 
a = 8'd247; b = 8'd247;  #10 
a = 8'd247; b = 8'd248;  #10 
a = 8'd247; b = 8'd249;  #10 
a = 8'd247; b = 8'd250;  #10 
a = 8'd247; b = 8'd251;  #10 
a = 8'd247; b = 8'd252;  #10 
a = 8'd247; b = 8'd253;  #10 
a = 8'd247; b = 8'd254;  #10 
a = 8'd247; b = 8'd255;  #10 
a = 8'd248; b = 8'd0;  #10 
a = 8'd248; b = 8'd1;  #10 
a = 8'd248; b = 8'd2;  #10 
a = 8'd248; b = 8'd3;  #10 
a = 8'd248; b = 8'd4;  #10 
a = 8'd248; b = 8'd5;  #10 
a = 8'd248; b = 8'd6;  #10 
a = 8'd248; b = 8'd7;  #10 
a = 8'd248; b = 8'd8;  #10 
a = 8'd248; b = 8'd9;  #10 
a = 8'd248; b = 8'd10;  #10 
a = 8'd248; b = 8'd11;  #10 
a = 8'd248; b = 8'd12;  #10 
a = 8'd248; b = 8'd13;  #10 
a = 8'd248; b = 8'd14;  #10 
a = 8'd248; b = 8'd15;  #10 
a = 8'd248; b = 8'd16;  #10 
a = 8'd248; b = 8'd17;  #10 
a = 8'd248; b = 8'd18;  #10 
a = 8'd248; b = 8'd19;  #10 
a = 8'd248; b = 8'd20;  #10 
a = 8'd248; b = 8'd21;  #10 
a = 8'd248; b = 8'd22;  #10 
a = 8'd248; b = 8'd23;  #10 
a = 8'd248; b = 8'd24;  #10 
a = 8'd248; b = 8'd25;  #10 
a = 8'd248; b = 8'd26;  #10 
a = 8'd248; b = 8'd27;  #10 
a = 8'd248; b = 8'd28;  #10 
a = 8'd248; b = 8'd29;  #10 
a = 8'd248; b = 8'd30;  #10 
a = 8'd248; b = 8'd31;  #10 
a = 8'd248; b = 8'd32;  #10 
a = 8'd248; b = 8'd33;  #10 
a = 8'd248; b = 8'd34;  #10 
a = 8'd248; b = 8'd35;  #10 
a = 8'd248; b = 8'd36;  #10 
a = 8'd248; b = 8'd37;  #10 
a = 8'd248; b = 8'd38;  #10 
a = 8'd248; b = 8'd39;  #10 
a = 8'd248; b = 8'd40;  #10 
a = 8'd248; b = 8'd41;  #10 
a = 8'd248; b = 8'd42;  #10 
a = 8'd248; b = 8'd43;  #10 
a = 8'd248; b = 8'd44;  #10 
a = 8'd248; b = 8'd45;  #10 
a = 8'd248; b = 8'd46;  #10 
a = 8'd248; b = 8'd47;  #10 
a = 8'd248; b = 8'd48;  #10 
a = 8'd248; b = 8'd49;  #10 
a = 8'd248; b = 8'd50;  #10 
a = 8'd248; b = 8'd51;  #10 
a = 8'd248; b = 8'd52;  #10 
a = 8'd248; b = 8'd53;  #10 
a = 8'd248; b = 8'd54;  #10 
a = 8'd248; b = 8'd55;  #10 
a = 8'd248; b = 8'd56;  #10 
a = 8'd248; b = 8'd57;  #10 
a = 8'd248; b = 8'd58;  #10 
a = 8'd248; b = 8'd59;  #10 
a = 8'd248; b = 8'd60;  #10 
a = 8'd248; b = 8'd61;  #10 
a = 8'd248; b = 8'd62;  #10 
a = 8'd248; b = 8'd63;  #10 
a = 8'd248; b = 8'd64;  #10 
a = 8'd248; b = 8'd65;  #10 
a = 8'd248; b = 8'd66;  #10 
a = 8'd248; b = 8'd67;  #10 
a = 8'd248; b = 8'd68;  #10 
a = 8'd248; b = 8'd69;  #10 
a = 8'd248; b = 8'd70;  #10 
a = 8'd248; b = 8'd71;  #10 
a = 8'd248; b = 8'd72;  #10 
a = 8'd248; b = 8'd73;  #10 
a = 8'd248; b = 8'd74;  #10 
a = 8'd248; b = 8'd75;  #10 
a = 8'd248; b = 8'd76;  #10 
a = 8'd248; b = 8'd77;  #10 
a = 8'd248; b = 8'd78;  #10 
a = 8'd248; b = 8'd79;  #10 
a = 8'd248; b = 8'd80;  #10 
a = 8'd248; b = 8'd81;  #10 
a = 8'd248; b = 8'd82;  #10 
a = 8'd248; b = 8'd83;  #10 
a = 8'd248; b = 8'd84;  #10 
a = 8'd248; b = 8'd85;  #10 
a = 8'd248; b = 8'd86;  #10 
a = 8'd248; b = 8'd87;  #10 
a = 8'd248; b = 8'd88;  #10 
a = 8'd248; b = 8'd89;  #10 
a = 8'd248; b = 8'd90;  #10 
a = 8'd248; b = 8'd91;  #10 
a = 8'd248; b = 8'd92;  #10 
a = 8'd248; b = 8'd93;  #10 
a = 8'd248; b = 8'd94;  #10 
a = 8'd248; b = 8'd95;  #10 
a = 8'd248; b = 8'd96;  #10 
a = 8'd248; b = 8'd97;  #10 
a = 8'd248; b = 8'd98;  #10 
a = 8'd248; b = 8'd99;  #10 
a = 8'd248; b = 8'd100;  #10 
a = 8'd248; b = 8'd101;  #10 
a = 8'd248; b = 8'd102;  #10 
a = 8'd248; b = 8'd103;  #10 
a = 8'd248; b = 8'd104;  #10 
a = 8'd248; b = 8'd105;  #10 
a = 8'd248; b = 8'd106;  #10 
a = 8'd248; b = 8'd107;  #10 
a = 8'd248; b = 8'd108;  #10 
a = 8'd248; b = 8'd109;  #10 
a = 8'd248; b = 8'd110;  #10 
a = 8'd248; b = 8'd111;  #10 
a = 8'd248; b = 8'd112;  #10 
a = 8'd248; b = 8'd113;  #10 
a = 8'd248; b = 8'd114;  #10 
a = 8'd248; b = 8'd115;  #10 
a = 8'd248; b = 8'd116;  #10 
a = 8'd248; b = 8'd117;  #10 
a = 8'd248; b = 8'd118;  #10 
a = 8'd248; b = 8'd119;  #10 
a = 8'd248; b = 8'd120;  #10 
a = 8'd248; b = 8'd121;  #10 
a = 8'd248; b = 8'd122;  #10 
a = 8'd248; b = 8'd123;  #10 
a = 8'd248; b = 8'd124;  #10 
a = 8'd248; b = 8'd125;  #10 
a = 8'd248; b = 8'd126;  #10 
a = 8'd248; b = 8'd127;  #10 
a = 8'd248; b = 8'd128;  #10 
a = 8'd248; b = 8'd129;  #10 
a = 8'd248; b = 8'd130;  #10 
a = 8'd248; b = 8'd131;  #10 
a = 8'd248; b = 8'd132;  #10 
a = 8'd248; b = 8'd133;  #10 
a = 8'd248; b = 8'd134;  #10 
a = 8'd248; b = 8'd135;  #10 
a = 8'd248; b = 8'd136;  #10 
a = 8'd248; b = 8'd137;  #10 
a = 8'd248; b = 8'd138;  #10 
a = 8'd248; b = 8'd139;  #10 
a = 8'd248; b = 8'd140;  #10 
a = 8'd248; b = 8'd141;  #10 
a = 8'd248; b = 8'd142;  #10 
a = 8'd248; b = 8'd143;  #10 
a = 8'd248; b = 8'd144;  #10 
a = 8'd248; b = 8'd145;  #10 
a = 8'd248; b = 8'd146;  #10 
a = 8'd248; b = 8'd147;  #10 
a = 8'd248; b = 8'd148;  #10 
a = 8'd248; b = 8'd149;  #10 
a = 8'd248; b = 8'd150;  #10 
a = 8'd248; b = 8'd151;  #10 
a = 8'd248; b = 8'd152;  #10 
a = 8'd248; b = 8'd153;  #10 
a = 8'd248; b = 8'd154;  #10 
a = 8'd248; b = 8'd155;  #10 
a = 8'd248; b = 8'd156;  #10 
a = 8'd248; b = 8'd157;  #10 
a = 8'd248; b = 8'd158;  #10 
a = 8'd248; b = 8'd159;  #10 
a = 8'd248; b = 8'd160;  #10 
a = 8'd248; b = 8'd161;  #10 
a = 8'd248; b = 8'd162;  #10 
a = 8'd248; b = 8'd163;  #10 
a = 8'd248; b = 8'd164;  #10 
a = 8'd248; b = 8'd165;  #10 
a = 8'd248; b = 8'd166;  #10 
a = 8'd248; b = 8'd167;  #10 
a = 8'd248; b = 8'd168;  #10 
a = 8'd248; b = 8'd169;  #10 
a = 8'd248; b = 8'd170;  #10 
a = 8'd248; b = 8'd171;  #10 
a = 8'd248; b = 8'd172;  #10 
a = 8'd248; b = 8'd173;  #10 
a = 8'd248; b = 8'd174;  #10 
a = 8'd248; b = 8'd175;  #10 
a = 8'd248; b = 8'd176;  #10 
a = 8'd248; b = 8'd177;  #10 
a = 8'd248; b = 8'd178;  #10 
a = 8'd248; b = 8'd179;  #10 
a = 8'd248; b = 8'd180;  #10 
a = 8'd248; b = 8'd181;  #10 
a = 8'd248; b = 8'd182;  #10 
a = 8'd248; b = 8'd183;  #10 
a = 8'd248; b = 8'd184;  #10 
a = 8'd248; b = 8'd185;  #10 
a = 8'd248; b = 8'd186;  #10 
a = 8'd248; b = 8'd187;  #10 
a = 8'd248; b = 8'd188;  #10 
a = 8'd248; b = 8'd189;  #10 
a = 8'd248; b = 8'd190;  #10 
a = 8'd248; b = 8'd191;  #10 
a = 8'd248; b = 8'd192;  #10 
a = 8'd248; b = 8'd193;  #10 
a = 8'd248; b = 8'd194;  #10 
a = 8'd248; b = 8'd195;  #10 
a = 8'd248; b = 8'd196;  #10 
a = 8'd248; b = 8'd197;  #10 
a = 8'd248; b = 8'd198;  #10 
a = 8'd248; b = 8'd199;  #10 
a = 8'd248; b = 8'd200;  #10 
a = 8'd248; b = 8'd201;  #10 
a = 8'd248; b = 8'd202;  #10 
a = 8'd248; b = 8'd203;  #10 
a = 8'd248; b = 8'd204;  #10 
a = 8'd248; b = 8'd205;  #10 
a = 8'd248; b = 8'd206;  #10 
a = 8'd248; b = 8'd207;  #10 
a = 8'd248; b = 8'd208;  #10 
a = 8'd248; b = 8'd209;  #10 
a = 8'd248; b = 8'd210;  #10 
a = 8'd248; b = 8'd211;  #10 
a = 8'd248; b = 8'd212;  #10 
a = 8'd248; b = 8'd213;  #10 
a = 8'd248; b = 8'd214;  #10 
a = 8'd248; b = 8'd215;  #10 
a = 8'd248; b = 8'd216;  #10 
a = 8'd248; b = 8'd217;  #10 
a = 8'd248; b = 8'd218;  #10 
a = 8'd248; b = 8'd219;  #10 
a = 8'd248; b = 8'd220;  #10 
a = 8'd248; b = 8'd221;  #10 
a = 8'd248; b = 8'd222;  #10 
a = 8'd248; b = 8'd223;  #10 
a = 8'd248; b = 8'd224;  #10 
a = 8'd248; b = 8'd225;  #10 
a = 8'd248; b = 8'd226;  #10 
a = 8'd248; b = 8'd227;  #10 
a = 8'd248; b = 8'd228;  #10 
a = 8'd248; b = 8'd229;  #10 
a = 8'd248; b = 8'd230;  #10 
a = 8'd248; b = 8'd231;  #10 
a = 8'd248; b = 8'd232;  #10 
a = 8'd248; b = 8'd233;  #10 
a = 8'd248; b = 8'd234;  #10 
a = 8'd248; b = 8'd235;  #10 
a = 8'd248; b = 8'd236;  #10 
a = 8'd248; b = 8'd237;  #10 
a = 8'd248; b = 8'd238;  #10 
a = 8'd248; b = 8'd239;  #10 
a = 8'd248; b = 8'd240;  #10 
a = 8'd248; b = 8'd241;  #10 
a = 8'd248; b = 8'd242;  #10 
a = 8'd248; b = 8'd243;  #10 
a = 8'd248; b = 8'd244;  #10 
a = 8'd248; b = 8'd245;  #10 
a = 8'd248; b = 8'd246;  #10 
a = 8'd248; b = 8'd247;  #10 
a = 8'd248; b = 8'd248;  #10 
a = 8'd248; b = 8'd249;  #10 
a = 8'd248; b = 8'd250;  #10 
a = 8'd248; b = 8'd251;  #10 
a = 8'd248; b = 8'd252;  #10 
a = 8'd248; b = 8'd253;  #10 
a = 8'd248; b = 8'd254;  #10 
a = 8'd248; b = 8'd255;  #10 
a = 8'd249; b = 8'd0;  #10 
a = 8'd249; b = 8'd1;  #10 
a = 8'd249; b = 8'd2;  #10 
a = 8'd249; b = 8'd3;  #10 
a = 8'd249; b = 8'd4;  #10 
a = 8'd249; b = 8'd5;  #10 
a = 8'd249; b = 8'd6;  #10 
a = 8'd249; b = 8'd7;  #10 
a = 8'd249; b = 8'd8;  #10 
a = 8'd249; b = 8'd9;  #10 
a = 8'd249; b = 8'd10;  #10 
a = 8'd249; b = 8'd11;  #10 
a = 8'd249; b = 8'd12;  #10 
a = 8'd249; b = 8'd13;  #10 
a = 8'd249; b = 8'd14;  #10 
a = 8'd249; b = 8'd15;  #10 
a = 8'd249; b = 8'd16;  #10 
a = 8'd249; b = 8'd17;  #10 
a = 8'd249; b = 8'd18;  #10 
a = 8'd249; b = 8'd19;  #10 
a = 8'd249; b = 8'd20;  #10 
a = 8'd249; b = 8'd21;  #10 
a = 8'd249; b = 8'd22;  #10 
a = 8'd249; b = 8'd23;  #10 
a = 8'd249; b = 8'd24;  #10 
a = 8'd249; b = 8'd25;  #10 
a = 8'd249; b = 8'd26;  #10 
a = 8'd249; b = 8'd27;  #10 
a = 8'd249; b = 8'd28;  #10 
a = 8'd249; b = 8'd29;  #10 
a = 8'd249; b = 8'd30;  #10 
a = 8'd249; b = 8'd31;  #10 
a = 8'd249; b = 8'd32;  #10 
a = 8'd249; b = 8'd33;  #10 
a = 8'd249; b = 8'd34;  #10 
a = 8'd249; b = 8'd35;  #10 
a = 8'd249; b = 8'd36;  #10 
a = 8'd249; b = 8'd37;  #10 
a = 8'd249; b = 8'd38;  #10 
a = 8'd249; b = 8'd39;  #10 
a = 8'd249; b = 8'd40;  #10 
a = 8'd249; b = 8'd41;  #10 
a = 8'd249; b = 8'd42;  #10 
a = 8'd249; b = 8'd43;  #10 
a = 8'd249; b = 8'd44;  #10 
a = 8'd249; b = 8'd45;  #10 
a = 8'd249; b = 8'd46;  #10 
a = 8'd249; b = 8'd47;  #10 
a = 8'd249; b = 8'd48;  #10 
a = 8'd249; b = 8'd49;  #10 
a = 8'd249; b = 8'd50;  #10 
a = 8'd249; b = 8'd51;  #10 
a = 8'd249; b = 8'd52;  #10 
a = 8'd249; b = 8'd53;  #10 
a = 8'd249; b = 8'd54;  #10 
a = 8'd249; b = 8'd55;  #10 
a = 8'd249; b = 8'd56;  #10 
a = 8'd249; b = 8'd57;  #10 
a = 8'd249; b = 8'd58;  #10 
a = 8'd249; b = 8'd59;  #10 
a = 8'd249; b = 8'd60;  #10 
a = 8'd249; b = 8'd61;  #10 
a = 8'd249; b = 8'd62;  #10 
a = 8'd249; b = 8'd63;  #10 
a = 8'd249; b = 8'd64;  #10 
a = 8'd249; b = 8'd65;  #10 
a = 8'd249; b = 8'd66;  #10 
a = 8'd249; b = 8'd67;  #10 
a = 8'd249; b = 8'd68;  #10 
a = 8'd249; b = 8'd69;  #10 
a = 8'd249; b = 8'd70;  #10 
a = 8'd249; b = 8'd71;  #10 
a = 8'd249; b = 8'd72;  #10 
a = 8'd249; b = 8'd73;  #10 
a = 8'd249; b = 8'd74;  #10 
a = 8'd249; b = 8'd75;  #10 
a = 8'd249; b = 8'd76;  #10 
a = 8'd249; b = 8'd77;  #10 
a = 8'd249; b = 8'd78;  #10 
a = 8'd249; b = 8'd79;  #10 
a = 8'd249; b = 8'd80;  #10 
a = 8'd249; b = 8'd81;  #10 
a = 8'd249; b = 8'd82;  #10 
a = 8'd249; b = 8'd83;  #10 
a = 8'd249; b = 8'd84;  #10 
a = 8'd249; b = 8'd85;  #10 
a = 8'd249; b = 8'd86;  #10 
a = 8'd249; b = 8'd87;  #10 
a = 8'd249; b = 8'd88;  #10 
a = 8'd249; b = 8'd89;  #10 
a = 8'd249; b = 8'd90;  #10 
a = 8'd249; b = 8'd91;  #10 
a = 8'd249; b = 8'd92;  #10 
a = 8'd249; b = 8'd93;  #10 
a = 8'd249; b = 8'd94;  #10 
a = 8'd249; b = 8'd95;  #10 
a = 8'd249; b = 8'd96;  #10 
a = 8'd249; b = 8'd97;  #10 
a = 8'd249; b = 8'd98;  #10 
a = 8'd249; b = 8'd99;  #10 
a = 8'd249; b = 8'd100;  #10 
a = 8'd249; b = 8'd101;  #10 
a = 8'd249; b = 8'd102;  #10 
a = 8'd249; b = 8'd103;  #10 
a = 8'd249; b = 8'd104;  #10 
a = 8'd249; b = 8'd105;  #10 
a = 8'd249; b = 8'd106;  #10 
a = 8'd249; b = 8'd107;  #10 
a = 8'd249; b = 8'd108;  #10 
a = 8'd249; b = 8'd109;  #10 
a = 8'd249; b = 8'd110;  #10 
a = 8'd249; b = 8'd111;  #10 
a = 8'd249; b = 8'd112;  #10 
a = 8'd249; b = 8'd113;  #10 
a = 8'd249; b = 8'd114;  #10 
a = 8'd249; b = 8'd115;  #10 
a = 8'd249; b = 8'd116;  #10 
a = 8'd249; b = 8'd117;  #10 
a = 8'd249; b = 8'd118;  #10 
a = 8'd249; b = 8'd119;  #10 
a = 8'd249; b = 8'd120;  #10 
a = 8'd249; b = 8'd121;  #10 
a = 8'd249; b = 8'd122;  #10 
a = 8'd249; b = 8'd123;  #10 
a = 8'd249; b = 8'd124;  #10 
a = 8'd249; b = 8'd125;  #10 
a = 8'd249; b = 8'd126;  #10 
a = 8'd249; b = 8'd127;  #10 
a = 8'd249; b = 8'd128;  #10 
a = 8'd249; b = 8'd129;  #10 
a = 8'd249; b = 8'd130;  #10 
a = 8'd249; b = 8'd131;  #10 
a = 8'd249; b = 8'd132;  #10 
a = 8'd249; b = 8'd133;  #10 
a = 8'd249; b = 8'd134;  #10 
a = 8'd249; b = 8'd135;  #10 
a = 8'd249; b = 8'd136;  #10 
a = 8'd249; b = 8'd137;  #10 
a = 8'd249; b = 8'd138;  #10 
a = 8'd249; b = 8'd139;  #10 
a = 8'd249; b = 8'd140;  #10 
a = 8'd249; b = 8'd141;  #10 
a = 8'd249; b = 8'd142;  #10 
a = 8'd249; b = 8'd143;  #10 
a = 8'd249; b = 8'd144;  #10 
a = 8'd249; b = 8'd145;  #10 
a = 8'd249; b = 8'd146;  #10 
a = 8'd249; b = 8'd147;  #10 
a = 8'd249; b = 8'd148;  #10 
a = 8'd249; b = 8'd149;  #10 
a = 8'd249; b = 8'd150;  #10 
a = 8'd249; b = 8'd151;  #10 
a = 8'd249; b = 8'd152;  #10 
a = 8'd249; b = 8'd153;  #10 
a = 8'd249; b = 8'd154;  #10 
a = 8'd249; b = 8'd155;  #10 
a = 8'd249; b = 8'd156;  #10 
a = 8'd249; b = 8'd157;  #10 
a = 8'd249; b = 8'd158;  #10 
a = 8'd249; b = 8'd159;  #10 
a = 8'd249; b = 8'd160;  #10 
a = 8'd249; b = 8'd161;  #10 
a = 8'd249; b = 8'd162;  #10 
a = 8'd249; b = 8'd163;  #10 
a = 8'd249; b = 8'd164;  #10 
a = 8'd249; b = 8'd165;  #10 
a = 8'd249; b = 8'd166;  #10 
a = 8'd249; b = 8'd167;  #10 
a = 8'd249; b = 8'd168;  #10 
a = 8'd249; b = 8'd169;  #10 
a = 8'd249; b = 8'd170;  #10 
a = 8'd249; b = 8'd171;  #10 
a = 8'd249; b = 8'd172;  #10 
a = 8'd249; b = 8'd173;  #10 
a = 8'd249; b = 8'd174;  #10 
a = 8'd249; b = 8'd175;  #10 
a = 8'd249; b = 8'd176;  #10 
a = 8'd249; b = 8'd177;  #10 
a = 8'd249; b = 8'd178;  #10 
a = 8'd249; b = 8'd179;  #10 
a = 8'd249; b = 8'd180;  #10 
a = 8'd249; b = 8'd181;  #10 
a = 8'd249; b = 8'd182;  #10 
a = 8'd249; b = 8'd183;  #10 
a = 8'd249; b = 8'd184;  #10 
a = 8'd249; b = 8'd185;  #10 
a = 8'd249; b = 8'd186;  #10 
a = 8'd249; b = 8'd187;  #10 
a = 8'd249; b = 8'd188;  #10 
a = 8'd249; b = 8'd189;  #10 
a = 8'd249; b = 8'd190;  #10 
a = 8'd249; b = 8'd191;  #10 
a = 8'd249; b = 8'd192;  #10 
a = 8'd249; b = 8'd193;  #10 
a = 8'd249; b = 8'd194;  #10 
a = 8'd249; b = 8'd195;  #10 
a = 8'd249; b = 8'd196;  #10 
a = 8'd249; b = 8'd197;  #10 
a = 8'd249; b = 8'd198;  #10 
a = 8'd249; b = 8'd199;  #10 
a = 8'd249; b = 8'd200;  #10 
a = 8'd249; b = 8'd201;  #10 
a = 8'd249; b = 8'd202;  #10 
a = 8'd249; b = 8'd203;  #10 
a = 8'd249; b = 8'd204;  #10 
a = 8'd249; b = 8'd205;  #10 
a = 8'd249; b = 8'd206;  #10 
a = 8'd249; b = 8'd207;  #10 
a = 8'd249; b = 8'd208;  #10 
a = 8'd249; b = 8'd209;  #10 
a = 8'd249; b = 8'd210;  #10 
a = 8'd249; b = 8'd211;  #10 
a = 8'd249; b = 8'd212;  #10 
a = 8'd249; b = 8'd213;  #10 
a = 8'd249; b = 8'd214;  #10 
a = 8'd249; b = 8'd215;  #10 
a = 8'd249; b = 8'd216;  #10 
a = 8'd249; b = 8'd217;  #10 
a = 8'd249; b = 8'd218;  #10 
a = 8'd249; b = 8'd219;  #10 
a = 8'd249; b = 8'd220;  #10 
a = 8'd249; b = 8'd221;  #10 
a = 8'd249; b = 8'd222;  #10 
a = 8'd249; b = 8'd223;  #10 
a = 8'd249; b = 8'd224;  #10 
a = 8'd249; b = 8'd225;  #10 
a = 8'd249; b = 8'd226;  #10 
a = 8'd249; b = 8'd227;  #10 
a = 8'd249; b = 8'd228;  #10 
a = 8'd249; b = 8'd229;  #10 
a = 8'd249; b = 8'd230;  #10 
a = 8'd249; b = 8'd231;  #10 
a = 8'd249; b = 8'd232;  #10 
a = 8'd249; b = 8'd233;  #10 
a = 8'd249; b = 8'd234;  #10 
a = 8'd249; b = 8'd235;  #10 
a = 8'd249; b = 8'd236;  #10 
a = 8'd249; b = 8'd237;  #10 
a = 8'd249; b = 8'd238;  #10 
a = 8'd249; b = 8'd239;  #10 
a = 8'd249; b = 8'd240;  #10 
a = 8'd249; b = 8'd241;  #10 
a = 8'd249; b = 8'd242;  #10 
a = 8'd249; b = 8'd243;  #10 
a = 8'd249; b = 8'd244;  #10 
a = 8'd249; b = 8'd245;  #10 
a = 8'd249; b = 8'd246;  #10 
a = 8'd249; b = 8'd247;  #10 
a = 8'd249; b = 8'd248;  #10 
a = 8'd249; b = 8'd249;  #10 
a = 8'd249; b = 8'd250;  #10 
a = 8'd249; b = 8'd251;  #10 
a = 8'd249; b = 8'd252;  #10 
a = 8'd249; b = 8'd253;  #10 
a = 8'd249; b = 8'd254;  #10 
a = 8'd249; b = 8'd255;  #10 
a = 8'd250; b = 8'd0;  #10 
a = 8'd250; b = 8'd1;  #10 
a = 8'd250; b = 8'd2;  #10 
a = 8'd250; b = 8'd3;  #10 
a = 8'd250; b = 8'd4;  #10 
a = 8'd250; b = 8'd5;  #10 
a = 8'd250; b = 8'd6;  #10 
a = 8'd250; b = 8'd7;  #10 
a = 8'd250; b = 8'd8;  #10 
a = 8'd250; b = 8'd9;  #10 
a = 8'd250; b = 8'd10;  #10 
a = 8'd250; b = 8'd11;  #10 
a = 8'd250; b = 8'd12;  #10 
a = 8'd250; b = 8'd13;  #10 
a = 8'd250; b = 8'd14;  #10 
a = 8'd250; b = 8'd15;  #10 
a = 8'd250; b = 8'd16;  #10 
a = 8'd250; b = 8'd17;  #10 
a = 8'd250; b = 8'd18;  #10 
a = 8'd250; b = 8'd19;  #10 
a = 8'd250; b = 8'd20;  #10 
a = 8'd250; b = 8'd21;  #10 
a = 8'd250; b = 8'd22;  #10 
a = 8'd250; b = 8'd23;  #10 
a = 8'd250; b = 8'd24;  #10 
a = 8'd250; b = 8'd25;  #10 
a = 8'd250; b = 8'd26;  #10 
a = 8'd250; b = 8'd27;  #10 
a = 8'd250; b = 8'd28;  #10 
a = 8'd250; b = 8'd29;  #10 
a = 8'd250; b = 8'd30;  #10 
a = 8'd250; b = 8'd31;  #10 
a = 8'd250; b = 8'd32;  #10 
a = 8'd250; b = 8'd33;  #10 
a = 8'd250; b = 8'd34;  #10 
a = 8'd250; b = 8'd35;  #10 
a = 8'd250; b = 8'd36;  #10 
a = 8'd250; b = 8'd37;  #10 
a = 8'd250; b = 8'd38;  #10 
a = 8'd250; b = 8'd39;  #10 
a = 8'd250; b = 8'd40;  #10 
a = 8'd250; b = 8'd41;  #10 
a = 8'd250; b = 8'd42;  #10 
a = 8'd250; b = 8'd43;  #10 
a = 8'd250; b = 8'd44;  #10 
a = 8'd250; b = 8'd45;  #10 
a = 8'd250; b = 8'd46;  #10 
a = 8'd250; b = 8'd47;  #10 
a = 8'd250; b = 8'd48;  #10 
a = 8'd250; b = 8'd49;  #10 
a = 8'd250; b = 8'd50;  #10 
a = 8'd250; b = 8'd51;  #10 
a = 8'd250; b = 8'd52;  #10 
a = 8'd250; b = 8'd53;  #10 
a = 8'd250; b = 8'd54;  #10 
a = 8'd250; b = 8'd55;  #10 
a = 8'd250; b = 8'd56;  #10 
a = 8'd250; b = 8'd57;  #10 
a = 8'd250; b = 8'd58;  #10 
a = 8'd250; b = 8'd59;  #10 
a = 8'd250; b = 8'd60;  #10 
a = 8'd250; b = 8'd61;  #10 
a = 8'd250; b = 8'd62;  #10 
a = 8'd250; b = 8'd63;  #10 
a = 8'd250; b = 8'd64;  #10 
a = 8'd250; b = 8'd65;  #10 
a = 8'd250; b = 8'd66;  #10 
a = 8'd250; b = 8'd67;  #10 
a = 8'd250; b = 8'd68;  #10 
a = 8'd250; b = 8'd69;  #10 
a = 8'd250; b = 8'd70;  #10 
a = 8'd250; b = 8'd71;  #10 
a = 8'd250; b = 8'd72;  #10 
a = 8'd250; b = 8'd73;  #10 
a = 8'd250; b = 8'd74;  #10 
a = 8'd250; b = 8'd75;  #10 
a = 8'd250; b = 8'd76;  #10 
a = 8'd250; b = 8'd77;  #10 
a = 8'd250; b = 8'd78;  #10 
a = 8'd250; b = 8'd79;  #10 
a = 8'd250; b = 8'd80;  #10 
a = 8'd250; b = 8'd81;  #10 
a = 8'd250; b = 8'd82;  #10 
a = 8'd250; b = 8'd83;  #10 
a = 8'd250; b = 8'd84;  #10 
a = 8'd250; b = 8'd85;  #10 
a = 8'd250; b = 8'd86;  #10 
a = 8'd250; b = 8'd87;  #10 
a = 8'd250; b = 8'd88;  #10 
a = 8'd250; b = 8'd89;  #10 
a = 8'd250; b = 8'd90;  #10 
a = 8'd250; b = 8'd91;  #10 
a = 8'd250; b = 8'd92;  #10 
a = 8'd250; b = 8'd93;  #10 
a = 8'd250; b = 8'd94;  #10 
a = 8'd250; b = 8'd95;  #10 
a = 8'd250; b = 8'd96;  #10 
a = 8'd250; b = 8'd97;  #10 
a = 8'd250; b = 8'd98;  #10 
a = 8'd250; b = 8'd99;  #10 
a = 8'd250; b = 8'd100;  #10 
a = 8'd250; b = 8'd101;  #10 
a = 8'd250; b = 8'd102;  #10 
a = 8'd250; b = 8'd103;  #10 
a = 8'd250; b = 8'd104;  #10 
a = 8'd250; b = 8'd105;  #10 
a = 8'd250; b = 8'd106;  #10 
a = 8'd250; b = 8'd107;  #10 
a = 8'd250; b = 8'd108;  #10 
a = 8'd250; b = 8'd109;  #10 
a = 8'd250; b = 8'd110;  #10 
a = 8'd250; b = 8'd111;  #10 
a = 8'd250; b = 8'd112;  #10 
a = 8'd250; b = 8'd113;  #10 
a = 8'd250; b = 8'd114;  #10 
a = 8'd250; b = 8'd115;  #10 
a = 8'd250; b = 8'd116;  #10 
a = 8'd250; b = 8'd117;  #10 
a = 8'd250; b = 8'd118;  #10 
a = 8'd250; b = 8'd119;  #10 
a = 8'd250; b = 8'd120;  #10 
a = 8'd250; b = 8'd121;  #10 
a = 8'd250; b = 8'd122;  #10 
a = 8'd250; b = 8'd123;  #10 
a = 8'd250; b = 8'd124;  #10 
a = 8'd250; b = 8'd125;  #10 
a = 8'd250; b = 8'd126;  #10 
a = 8'd250; b = 8'd127;  #10 
a = 8'd250; b = 8'd128;  #10 
a = 8'd250; b = 8'd129;  #10 
a = 8'd250; b = 8'd130;  #10 
a = 8'd250; b = 8'd131;  #10 
a = 8'd250; b = 8'd132;  #10 
a = 8'd250; b = 8'd133;  #10 
a = 8'd250; b = 8'd134;  #10 
a = 8'd250; b = 8'd135;  #10 
a = 8'd250; b = 8'd136;  #10 
a = 8'd250; b = 8'd137;  #10 
a = 8'd250; b = 8'd138;  #10 
a = 8'd250; b = 8'd139;  #10 
a = 8'd250; b = 8'd140;  #10 
a = 8'd250; b = 8'd141;  #10 
a = 8'd250; b = 8'd142;  #10 
a = 8'd250; b = 8'd143;  #10 
a = 8'd250; b = 8'd144;  #10 
a = 8'd250; b = 8'd145;  #10 
a = 8'd250; b = 8'd146;  #10 
a = 8'd250; b = 8'd147;  #10 
a = 8'd250; b = 8'd148;  #10 
a = 8'd250; b = 8'd149;  #10 
a = 8'd250; b = 8'd150;  #10 
a = 8'd250; b = 8'd151;  #10 
a = 8'd250; b = 8'd152;  #10 
a = 8'd250; b = 8'd153;  #10 
a = 8'd250; b = 8'd154;  #10 
a = 8'd250; b = 8'd155;  #10 
a = 8'd250; b = 8'd156;  #10 
a = 8'd250; b = 8'd157;  #10 
a = 8'd250; b = 8'd158;  #10 
a = 8'd250; b = 8'd159;  #10 
a = 8'd250; b = 8'd160;  #10 
a = 8'd250; b = 8'd161;  #10 
a = 8'd250; b = 8'd162;  #10 
a = 8'd250; b = 8'd163;  #10 
a = 8'd250; b = 8'd164;  #10 
a = 8'd250; b = 8'd165;  #10 
a = 8'd250; b = 8'd166;  #10 
a = 8'd250; b = 8'd167;  #10 
a = 8'd250; b = 8'd168;  #10 
a = 8'd250; b = 8'd169;  #10 
a = 8'd250; b = 8'd170;  #10 
a = 8'd250; b = 8'd171;  #10 
a = 8'd250; b = 8'd172;  #10 
a = 8'd250; b = 8'd173;  #10 
a = 8'd250; b = 8'd174;  #10 
a = 8'd250; b = 8'd175;  #10 
a = 8'd250; b = 8'd176;  #10 
a = 8'd250; b = 8'd177;  #10 
a = 8'd250; b = 8'd178;  #10 
a = 8'd250; b = 8'd179;  #10 
a = 8'd250; b = 8'd180;  #10 
a = 8'd250; b = 8'd181;  #10 
a = 8'd250; b = 8'd182;  #10 
a = 8'd250; b = 8'd183;  #10 
a = 8'd250; b = 8'd184;  #10 
a = 8'd250; b = 8'd185;  #10 
a = 8'd250; b = 8'd186;  #10 
a = 8'd250; b = 8'd187;  #10 
a = 8'd250; b = 8'd188;  #10 
a = 8'd250; b = 8'd189;  #10 
a = 8'd250; b = 8'd190;  #10 
a = 8'd250; b = 8'd191;  #10 
a = 8'd250; b = 8'd192;  #10 
a = 8'd250; b = 8'd193;  #10 
a = 8'd250; b = 8'd194;  #10 
a = 8'd250; b = 8'd195;  #10 
a = 8'd250; b = 8'd196;  #10 
a = 8'd250; b = 8'd197;  #10 
a = 8'd250; b = 8'd198;  #10 
a = 8'd250; b = 8'd199;  #10 
a = 8'd250; b = 8'd200;  #10 
a = 8'd250; b = 8'd201;  #10 
a = 8'd250; b = 8'd202;  #10 
a = 8'd250; b = 8'd203;  #10 
a = 8'd250; b = 8'd204;  #10 
a = 8'd250; b = 8'd205;  #10 
a = 8'd250; b = 8'd206;  #10 
a = 8'd250; b = 8'd207;  #10 
a = 8'd250; b = 8'd208;  #10 
a = 8'd250; b = 8'd209;  #10 
a = 8'd250; b = 8'd210;  #10 
a = 8'd250; b = 8'd211;  #10 
a = 8'd250; b = 8'd212;  #10 
a = 8'd250; b = 8'd213;  #10 
a = 8'd250; b = 8'd214;  #10 
a = 8'd250; b = 8'd215;  #10 
a = 8'd250; b = 8'd216;  #10 
a = 8'd250; b = 8'd217;  #10 
a = 8'd250; b = 8'd218;  #10 
a = 8'd250; b = 8'd219;  #10 
a = 8'd250; b = 8'd220;  #10 
a = 8'd250; b = 8'd221;  #10 
a = 8'd250; b = 8'd222;  #10 
a = 8'd250; b = 8'd223;  #10 
a = 8'd250; b = 8'd224;  #10 
a = 8'd250; b = 8'd225;  #10 
a = 8'd250; b = 8'd226;  #10 
a = 8'd250; b = 8'd227;  #10 
a = 8'd250; b = 8'd228;  #10 
a = 8'd250; b = 8'd229;  #10 
a = 8'd250; b = 8'd230;  #10 
a = 8'd250; b = 8'd231;  #10 
a = 8'd250; b = 8'd232;  #10 
a = 8'd250; b = 8'd233;  #10 
a = 8'd250; b = 8'd234;  #10 
a = 8'd250; b = 8'd235;  #10 
a = 8'd250; b = 8'd236;  #10 
a = 8'd250; b = 8'd237;  #10 
a = 8'd250; b = 8'd238;  #10 
a = 8'd250; b = 8'd239;  #10 
a = 8'd250; b = 8'd240;  #10 
a = 8'd250; b = 8'd241;  #10 
a = 8'd250; b = 8'd242;  #10 
a = 8'd250; b = 8'd243;  #10 
a = 8'd250; b = 8'd244;  #10 
a = 8'd250; b = 8'd245;  #10 
a = 8'd250; b = 8'd246;  #10 
a = 8'd250; b = 8'd247;  #10 
a = 8'd250; b = 8'd248;  #10 
a = 8'd250; b = 8'd249;  #10 
a = 8'd250; b = 8'd250;  #10 
a = 8'd250; b = 8'd251;  #10 
a = 8'd250; b = 8'd252;  #10 
a = 8'd250; b = 8'd253;  #10 
a = 8'd250; b = 8'd254;  #10 
a = 8'd250; b = 8'd255;  #10 
a = 8'd251; b = 8'd0;  #10 
a = 8'd251; b = 8'd1;  #10 
a = 8'd251; b = 8'd2;  #10 
a = 8'd251; b = 8'd3;  #10 
a = 8'd251; b = 8'd4;  #10 
a = 8'd251; b = 8'd5;  #10 
a = 8'd251; b = 8'd6;  #10 
a = 8'd251; b = 8'd7;  #10 
a = 8'd251; b = 8'd8;  #10 
a = 8'd251; b = 8'd9;  #10 
a = 8'd251; b = 8'd10;  #10 
a = 8'd251; b = 8'd11;  #10 
a = 8'd251; b = 8'd12;  #10 
a = 8'd251; b = 8'd13;  #10 
a = 8'd251; b = 8'd14;  #10 
a = 8'd251; b = 8'd15;  #10 
a = 8'd251; b = 8'd16;  #10 
a = 8'd251; b = 8'd17;  #10 
a = 8'd251; b = 8'd18;  #10 
a = 8'd251; b = 8'd19;  #10 
a = 8'd251; b = 8'd20;  #10 
a = 8'd251; b = 8'd21;  #10 
a = 8'd251; b = 8'd22;  #10 
a = 8'd251; b = 8'd23;  #10 
a = 8'd251; b = 8'd24;  #10 
a = 8'd251; b = 8'd25;  #10 
a = 8'd251; b = 8'd26;  #10 
a = 8'd251; b = 8'd27;  #10 
a = 8'd251; b = 8'd28;  #10 
a = 8'd251; b = 8'd29;  #10 
a = 8'd251; b = 8'd30;  #10 
a = 8'd251; b = 8'd31;  #10 
a = 8'd251; b = 8'd32;  #10 
a = 8'd251; b = 8'd33;  #10 
a = 8'd251; b = 8'd34;  #10 
a = 8'd251; b = 8'd35;  #10 
a = 8'd251; b = 8'd36;  #10 
a = 8'd251; b = 8'd37;  #10 
a = 8'd251; b = 8'd38;  #10 
a = 8'd251; b = 8'd39;  #10 
a = 8'd251; b = 8'd40;  #10 
a = 8'd251; b = 8'd41;  #10 
a = 8'd251; b = 8'd42;  #10 
a = 8'd251; b = 8'd43;  #10 
a = 8'd251; b = 8'd44;  #10 
a = 8'd251; b = 8'd45;  #10 
a = 8'd251; b = 8'd46;  #10 
a = 8'd251; b = 8'd47;  #10 
a = 8'd251; b = 8'd48;  #10 
a = 8'd251; b = 8'd49;  #10 
a = 8'd251; b = 8'd50;  #10 
a = 8'd251; b = 8'd51;  #10 
a = 8'd251; b = 8'd52;  #10 
a = 8'd251; b = 8'd53;  #10 
a = 8'd251; b = 8'd54;  #10 
a = 8'd251; b = 8'd55;  #10 
a = 8'd251; b = 8'd56;  #10 
a = 8'd251; b = 8'd57;  #10 
a = 8'd251; b = 8'd58;  #10 
a = 8'd251; b = 8'd59;  #10 
a = 8'd251; b = 8'd60;  #10 
a = 8'd251; b = 8'd61;  #10 
a = 8'd251; b = 8'd62;  #10 
a = 8'd251; b = 8'd63;  #10 
a = 8'd251; b = 8'd64;  #10 
a = 8'd251; b = 8'd65;  #10 
a = 8'd251; b = 8'd66;  #10 
a = 8'd251; b = 8'd67;  #10 
a = 8'd251; b = 8'd68;  #10 
a = 8'd251; b = 8'd69;  #10 
a = 8'd251; b = 8'd70;  #10 
a = 8'd251; b = 8'd71;  #10 
a = 8'd251; b = 8'd72;  #10 
a = 8'd251; b = 8'd73;  #10 
a = 8'd251; b = 8'd74;  #10 
a = 8'd251; b = 8'd75;  #10 
a = 8'd251; b = 8'd76;  #10 
a = 8'd251; b = 8'd77;  #10 
a = 8'd251; b = 8'd78;  #10 
a = 8'd251; b = 8'd79;  #10 
a = 8'd251; b = 8'd80;  #10 
a = 8'd251; b = 8'd81;  #10 
a = 8'd251; b = 8'd82;  #10 
a = 8'd251; b = 8'd83;  #10 
a = 8'd251; b = 8'd84;  #10 
a = 8'd251; b = 8'd85;  #10 
a = 8'd251; b = 8'd86;  #10 
a = 8'd251; b = 8'd87;  #10 
a = 8'd251; b = 8'd88;  #10 
a = 8'd251; b = 8'd89;  #10 
a = 8'd251; b = 8'd90;  #10 
a = 8'd251; b = 8'd91;  #10 
a = 8'd251; b = 8'd92;  #10 
a = 8'd251; b = 8'd93;  #10 
a = 8'd251; b = 8'd94;  #10 
a = 8'd251; b = 8'd95;  #10 
a = 8'd251; b = 8'd96;  #10 
a = 8'd251; b = 8'd97;  #10 
a = 8'd251; b = 8'd98;  #10 
a = 8'd251; b = 8'd99;  #10 
a = 8'd251; b = 8'd100;  #10 
a = 8'd251; b = 8'd101;  #10 
a = 8'd251; b = 8'd102;  #10 
a = 8'd251; b = 8'd103;  #10 
a = 8'd251; b = 8'd104;  #10 
a = 8'd251; b = 8'd105;  #10 
a = 8'd251; b = 8'd106;  #10 
a = 8'd251; b = 8'd107;  #10 
a = 8'd251; b = 8'd108;  #10 
a = 8'd251; b = 8'd109;  #10 
a = 8'd251; b = 8'd110;  #10 
a = 8'd251; b = 8'd111;  #10 
a = 8'd251; b = 8'd112;  #10 
a = 8'd251; b = 8'd113;  #10 
a = 8'd251; b = 8'd114;  #10 
a = 8'd251; b = 8'd115;  #10 
a = 8'd251; b = 8'd116;  #10 
a = 8'd251; b = 8'd117;  #10 
a = 8'd251; b = 8'd118;  #10 
a = 8'd251; b = 8'd119;  #10 
a = 8'd251; b = 8'd120;  #10 
a = 8'd251; b = 8'd121;  #10 
a = 8'd251; b = 8'd122;  #10 
a = 8'd251; b = 8'd123;  #10 
a = 8'd251; b = 8'd124;  #10 
a = 8'd251; b = 8'd125;  #10 
a = 8'd251; b = 8'd126;  #10 
a = 8'd251; b = 8'd127;  #10 
a = 8'd251; b = 8'd128;  #10 
a = 8'd251; b = 8'd129;  #10 
a = 8'd251; b = 8'd130;  #10 
a = 8'd251; b = 8'd131;  #10 
a = 8'd251; b = 8'd132;  #10 
a = 8'd251; b = 8'd133;  #10 
a = 8'd251; b = 8'd134;  #10 
a = 8'd251; b = 8'd135;  #10 
a = 8'd251; b = 8'd136;  #10 
a = 8'd251; b = 8'd137;  #10 
a = 8'd251; b = 8'd138;  #10 
a = 8'd251; b = 8'd139;  #10 
a = 8'd251; b = 8'd140;  #10 
a = 8'd251; b = 8'd141;  #10 
a = 8'd251; b = 8'd142;  #10 
a = 8'd251; b = 8'd143;  #10 
a = 8'd251; b = 8'd144;  #10 
a = 8'd251; b = 8'd145;  #10 
a = 8'd251; b = 8'd146;  #10 
a = 8'd251; b = 8'd147;  #10 
a = 8'd251; b = 8'd148;  #10 
a = 8'd251; b = 8'd149;  #10 
a = 8'd251; b = 8'd150;  #10 
a = 8'd251; b = 8'd151;  #10 
a = 8'd251; b = 8'd152;  #10 
a = 8'd251; b = 8'd153;  #10 
a = 8'd251; b = 8'd154;  #10 
a = 8'd251; b = 8'd155;  #10 
a = 8'd251; b = 8'd156;  #10 
a = 8'd251; b = 8'd157;  #10 
a = 8'd251; b = 8'd158;  #10 
a = 8'd251; b = 8'd159;  #10 
a = 8'd251; b = 8'd160;  #10 
a = 8'd251; b = 8'd161;  #10 
a = 8'd251; b = 8'd162;  #10 
a = 8'd251; b = 8'd163;  #10 
a = 8'd251; b = 8'd164;  #10 
a = 8'd251; b = 8'd165;  #10 
a = 8'd251; b = 8'd166;  #10 
a = 8'd251; b = 8'd167;  #10 
a = 8'd251; b = 8'd168;  #10 
a = 8'd251; b = 8'd169;  #10 
a = 8'd251; b = 8'd170;  #10 
a = 8'd251; b = 8'd171;  #10 
a = 8'd251; b = 8'd172;  #10 
a = 8'd251; b = 8'd173;  #10 
a = 8'd251; b = 8'd174;  #10 
a = 8'd251; b = 8'd175;  #10 
a = 8'd251; b = 8'd176;  #10 
a = 8'd251; b = 8'd177;  #10 
a = 8'd251; b = 8'd178;  #10 
a = 8'd251; b = 8'd179;  #10 
a = 8'd251; b = 8'd180;  #10 
a = 8'd251; b = 8'd181;  #10 
a = 8'd251; b = 8'd182;  #10 
a = 8'd251; b = 8'd183;  #10 
a = 8'd251; b = 8'd184;  #10 
a = 8'd251; b = 8'd185;  #10 
a = 8'd251; b = 8'd186;  #10 
a = 8'd251; b = 8'd187;  #10 
a = 8'd251; b = 8'd188;  #10 
a = 8'd251; b = 8'd189;  #10 
a = 8'd251; b = 8'd190;  #10 
a = 8'd251; b = 8'd191;  #10 
a = 8'd251; b = 8'd192;  #10 
a = 8'd251; b = 8'd193;  #10 
a = 8'd251; b = 8'd194;  #10 
a = 8'd251; b = 8'd195;  #10 
a = 8'd251; b = 8'd196;  #10 
a = 8'd251; b = 8'd197;  #10 
a = 8'd251; b = 8'd198;  #10 
a = 8'd251; b = 8'd199;  #10 
a = 8'd251; b = 8'd200;  #10 
a = 8'd251; b = 8'd201;  #10 
a = 8'd251; b = 8'd202;  #10 
a = 8'd251; b = 8'd203;  #10 
a = 8'd251; b = 8'd204;  #10 
a = 8'd251; b = 8'd205;  #10 
a = 8'd251; b = 8'd206;  #10 
a = 8'd251; b = 8'd207;  #10 
a = 8'd251; b = 8'd208;  #10 
a = 8'd251; b = 8'd209;  #10 
a = 8'd251; b = 8'd210;  #10 
a = 8'd251; b = 8'd211;  #10 
a = 8'd251; b = 8'd212;  #10 
a = 8'd251; b = 8'd213;  #10 
a = 8'd251; b = 8'd214;  #10 
a = 8'd251; b = 8'd215;  #10 
a = 8'd251; b = 8'd216;  #10 
a = 8'd251; b = 8'd217;  #10 
a = 8'd251; b = 8'd218;  #10 
a = 8'd251; b = 8'd219;  #10 
a = 8'd251; b = 8'd220;  #10 
a = 8'd251; b = 8'd221;  #10 
a = 8'd251; b = 8'd222;  #10 
a = 8'd251; b = 8'd223;  #10 
a = 8'd251; b = 8'd224;  #10 
a = 8'd251; b = 8'd225;  #10 
a = 8'd251; b = 8'd226;  #10 
a = 8'd251; b = 8'd227;  #10 
a = 8'd251; b = 8'd228;  #10 
a = 8'd251; b = 8'd229;  #10 
a = 8'd251; b = 8'd230;  #10 
a = 8'd251; b = 8'd231;  #10 
a = 8'd251; b = 8'd232;  #10 
a = 8'd251; b = 8'd233;  #10 
a = 8'd251; b = 8'd234;  #10 
a = 8'd251; b = 8'd235;  #10 
a = 8'd251; b = 8'd236;  #10 
a = 8'd251; b = 8'd237;  #10 
a = 8'd251; b = 8'd238;  #10 
a = 8'd251; b = 8'd239;  #10 
a = 8'd251; b = 8'd240;  #10 
a = 8'd251; b = 8'd241;  #10 
a = 8'd251; b = 8'd242;  #10 
a = 8'd251; b = 8'd243;  #10 
a = 8'd251; b = 8'd244;  #10 
a = 8'd251; b = 8'd245;  #10 
a = 8'd251; b = 8'd246;  #10 
a = 8'd251; b = 8'd247;  #10 
a = 8'd251; b = 8'd248;  #10 
a = 8'd251; b = 8'd249;  #10 
a = 8'd251; b = 8'd250;  #10 
a = 8'd251; b = 8'd251;  #10 
a = 8'd251; b = 8'd252;  #10 
a = 8'd251; b = 8'd253;  #10 
a = 8'd251; b = 8'd254;  #10 
a = 8'd251; b = 8'd255;  #10 
a = 8'd252; b = 8'd0;  #10 
a = 8'd252; b = 8'd1;  #10 
a = 8'd252; b = 8'd2;  #10 
a = 8'd252; b = 8'd3;  #10 
a = 8'd252; b = 8'd4;  #10 
a = 8'd252; b = 8'd5;  #10 
a = 8'd252; b = 8'd6;  #10 
a = 8'd252; b = 8'd7;  #10 
a = 8'd252; b = 8'd8;  #10 
a = 8'd252; b = 8'd9;  #10 
a = 8'd252; b = 8'd10;  #10 
a = 8'd252; b = 8'd11;  #10 
a = 8'd252; b = 8'd12;  #10 
a = 8'd252; b = 8'd13;  #10 
a = 8'd252; b = 8'd14;  #10 
a = 8'd252; b = 8'd15;  #10 
a = 8'd252; b = 8'd16;  #10 
a = 8'd252; b = 8'd17;  #10 
a = 8'd252; b = 8'd18;  #10 
a = 8'd252; b = 8'd19;  #10 
a = 8'd252; b = 8'd20;  #10 
a = 8'd252; b = 8'd21;  #10 
a = 8'd252; b = 8'd22;  #10 
a = 8'd252; b = 8'd23;  #10 
a = 8'd252; b = 8'd24;  #10 
a = 8'd252; b = 8'd25;  #10 
a = 8'd252; b = 8'd26;  #10 
a = 8'd252; b = 8'd27;  #10 
a = 8'd252; b = 8'd28;  #10 
a = 8'd252; b = 8'd29;  #10 
a = 8'd252; b = 8'd30;  #10 
a = 8'd252; b = 8'd31;  #10 
a = 8'd252; b = 8'd32;  #10 
a = 8'd252; b = 8'd33;  #10 
a = 8'd252; b = 8'd34;  #10 
a = 8'd252; b = 8'd35;  #10 
a = 8'd252; b = 8'd36;  #10 
a = 8'd252; b = 8'd37;  #10 
a = 8'd252; b = 8'd38;  #10 
a = 8'd252; b = 8'd39;  #10 
a = 8'd252; b = 8'd40;  #10 
a = 8'd252; b = 8'd41;  #10 
a = 8'd252; b = 8'd42;  #10 
a = 8'd252; b = 8'd43;  #10 
a = 8'd252; b = 8'd44;  #10 
a = 8'd252; b = 8'd45;  #10 
a = 8'd252; b = 8'd46;  #10 
a = 8'd252; b = 8'd47;  #10 
a = 8'd252; b = 8'd48;  #10 
a = 8'd252; b = 8'd49;  #10 
a = 8'd252; b = 8'd50;  #10 
a = 8'd252; b = 8'd51;  #10 
a = 8'd252; b = 8'd52;  #10 
a = 8'd252; b = 8'd53;  #10 
a = 8'd252; b = 8'd54;  #10 
a = 8'd252; b = 8'd55;  #10 
a = 8'd252; b = 8'd56;  #10 
a = 8'd252; b = 8'd57;  #10 
a = 8'd252; b = 8'd58;  #10 
a = 8'd252; b = 8'd59;  #10 
a = 8'd252; b = 8'd60;  #10 
a = 8'd252; b = 8'd61;  #10 
a = 8'd252; b = 8'd62;  #10 
a = 8'd252; b = 8'd63;  #10 
a = 8'd252; b = 8'd64;  #10 
a = 8'd252; b = 8'd65;  #10 
a = 8'd252; b = 8'd66;  #10 
a = 8'd252; b = 8'd67;  #10 
a = 8'd252; b = 8'd68;  #10 
a = 8'd252; b = 8'd69;  #10 
a = 8'd252; b = 8'd70;  #10 
a = 8'd252; b = 8'd71;  #10 
a = 8'd252; b = 8'd72;  #10 
a = 8'd252; b = 8'd73;  #10 
a = 8'd252; b = 8'd74;  #10 
a = 8'd252; b = 8'd75;  #10 
a = 8'd252; b = 8'd76;  #10 
a = 8'd252; b = 8'd77;  #10 
a = 8'd252; b = 8'd78;  #10 
a = 8'd252; b = 8'd79;  #10 
a = 8'd252; b = 8'd80;  #10 
a = 8'd252; b = 8'd81;  #10 
a = 8'd252; b = 8'd82;  #10 
a = 8'd252; b = 8'd83;  #10 
a = 8'd252; b = 8'd84;  #10 
a = 8'd252; b = 8'd85;  #10 
a = 8'd252; b = 8'd86;  #10 
a = 8'd252; b = 8'd87;  #10 
a = 8'd252; b = 8'd88;  #10 
a = 8'd252; b = 8'd89;  #10 
a = 8'd252; b = 8'd90;  #10 
a = 8'd252; b = 8'd91;  #10 
a = 8'd252; b = 8'd92;  #10 
a = 8'd252; b = 8'd93;  #10 
a = 8'd252; b = 8'd94;  #10 
a = 8'd252; b = 8'd95;  #10 
a = 8'd252; b = 8'd96;  #10 
a = 8'd252; b = 8'd97;  #10 
a = 8'd252; b = 8'd98;  #10 
a = 8'd252; b = 8'd99;  #10 
a = 8'd252; b = 8'd100;  #10 
a = 8'd252; b = 8'd101;  #10 
a = 8'd252; b = 8'd102;  #10 
a = 8'd252; b = 8'd103;  #10 
a = 8'd252; b = 8'd104;  #10 
a = 8'd252; b = 8'd105;  #10 
a = 8'd252; b = 8'd106;  #10 
a = 8'd252; b = 8'd107;  #10 
a = 8'd252; b = 8'd108;  #10 
a = 8'd252; b = 8'd109;  #10 
a = 8'd252; b = 8'd110;  #10 
a = 8'd252; b = 8'd111;  #10 
a = 8'd252; b = 8'd112;  #10 
a = 8'd252; b = 8'd113;  #10 
a = 8'd252; b = 8'd114;  #10 
a = 8'd252; b = 8'd115;  #10 
a = 8'd252; b = 8'd116;  #10 
a = 8'd252; b = 8'd117;  #10 
a = 8'd252; b = 8'd118;  #10 
a = 8'd252; b = 8'd119;  #10 
a = 8'd252; b = 8'd120;  #10 
a = 8'd252; b = 8'd121;  #10 
a = 8'd252; b = 8'd122;  #10 
a = 8'd252; b = 8'd123;  #10 
a = 8'd252; b = 8'd124;  #10 
a = 8'd252; b = 8'd125;  #10 
a = 8'd252; b = 8'd126;  #10 
a = 8'd252; b = 8'd127;  #10 
a = 8'd252; b = 8'd128;  #10 
a = 8'd252; b = 8'd129;  #10 
a = 8'd252; b = 8'd130;  #10 
a = 8'd252; b = 8'd131;  #10 
a = 8'd252; b = 8'd132;  #10 
a = 8'd252; b = 8'd133;  #10 
a = 8'd252; b = 8'd134;  #10 
a = 8'd252; b = 8'd135;  #10 
a = 8'd252; b = 8'd136;  #10 
a = 8'd252; b = 8'd137;  #10 
a = 8'd252; b = 8'd138;  #10 
a = 8'd252; b = 8'd139;  #10 
a = 8'd252; b = 8'd140;  #10 
a = 8'd252; b = 8'd141;  #10 
a = 8'd252; b = 8'd142;  #10 
a = 8'd252; b = 8'd143;  #10 
a = 8'd252; b = 8'd144;  #10 
a = 8'd252; b = 8'd145;  #10 
a = 8'd252; b = 8'd146;  #10 
a = 8'd252; b = 8'd147;  #10 
a = 8'd252; b = 8'd148;  #10 
a = 8'd252; b = 8'd149;  #10 
a = 8'd252; b = 8'd150;  #10 
a = 8'd252; b = 8'd151;  #10 
a = 8'd252; b = 8'd152;  #10 
a = 8'd252; b = 8'd153;  #10 
a = 8'd252; b = 8'd154;  #10 
a = 8'd252; b = 8'd155;  #10 
a = 8'd252; b = 8'd156;  #10 
a = 8'd252; b = 8'd157;  #10 
a = 8'd252; b = 8'd158;  #10 
a = 8'd252; b = 8'd159;  #10 
a = 8'd252; b = 8'd160;  #10 
a = 8'd252; b = 8'd161;  #10 
a = 8'd252; b = 8'd162;  #10 
a = 8'd252; b = 8'd163;  #10 
a = 8'd252; b = 8'd164;  #10 
a = 8'd252; b = 8'd165;  #10 
a = 8'd252; b = 8'd166;  #10 
a = 8'd252; b = 8'd167;  #10 
a = 8'd252; b = 8'd168;  #10 
a = 8'd252; b = 8'd169;  #10 
a = 8'd252; b = 8'd170;  #10 
a = 8'd252; b = 8'd171;  #10 
a = 8'd252; b = 8'd172;  #10 
a = 8'd252; b = 8'd173;  #10 
a = 8'd252; b = 8'd174;  #10 
a = 8'd252; b = 8'd175;  #10 
a = 8'd252; b = 8'd176;  #10 
a = 8'd252; b = 8'd177;  #10 
a = 8'd252; b = 8'd178;  #10 
a = 8'd252; b = 8'd179;  #10 
a = 8'd252; b = 8'd180;  #10 
a = 8'd252; b = 8'd181;  #10 
a = 8'd252; b = 8'd182;  #10 
a = 8'd252; b = 8'd183;  #10 
a = 8'd252; b = 8'd184;  #10 
a = 8'd252; b = 8'd185;  #10 
a = 8'd252; b = 8'd186;  #10 
a = 8'd252; b = 8'd187;  #10 
a = 8'd252; b = 8'd188;  #10 
a = 8'd252; b = 8'd189;  #10 
a = 8'd252; b = 8'd190;  #10 
a = 8'd252; b = 8'd191;  #10 
a = 8'd252; b = 8'd192;  #10 
a = 8'd252; b = 8'd193;  #10 
a = 8'd252; b = 8'd194;  #10 
a = 8'd252; b = 8'd195;  #10 
a = 8'd252; b = 8'd196;  #10 
a = 8'd252; b = 8'd197;  #10 
a = 8'd252; b = 8'd198;  #10 
a = 8'd252; b = 8'd199;  #10 
a = 8'd252; b = 8'd200;  #10 
a = 8'd252; b = 8'd201;  #10 
a = 8'd252; b = 8'd202;  #10 
a = 8'd252; b = 8'd203;  #10 
a = 8'd252; b = 8'd204;  #10 
a = 8'd252; b = 8'd205;  #10 
a = 8'd252; b = 8'd206;  #10 
a = 8'd252; b = 8'd207;  #10 
a = 8'd252; b = 8'd208;  #10 
a = 8'd252; b = 8'd209;  #10 
a = 8'd252; b = 8'd210;  #10 
a = 8'd252; b = 8'd211;  #10 
a = 8'd252; b = 8'd212;  #10 
a = 8'd252; b = 8'd213;  #10 
a = 8'd252; b = 8'd214;  #10 
a = 8'd252; b = 8'd215;  #10 
a = 8'd252; b = 8'd216;  #10 
a = 8'd252; b = 8'd217;  #10 
a = 8'd252; b = 8'd218;  #10 
a = 8'd252; b = 8'd219;  #10 
a = 8'd252; b = 8'd220;  #10 
a = 8'd252; b = 8'd221;  #10 
a = 8'd252; b = 8'd222;  #10 
a = 8'd252; b = 8'd223;  #10 
a = 8'd252; b = 8'd224;  #10 
a = 8'd252; b = 8'd225;  #10 
a = 8'd252; b = 8'd226;  #10 
a = 8'd252; b = 8'd227;  #10 
a = 8'd252; b = 8'd228;  #10 
a = 8'd252; b = 8'd229;  #10 
a = 8'd252; b = 8'd230;  #10 
a = 8'd252; b = 8'd231;  #10 
a = 8'd252; b = 8'd232;  #10 
a = 8'd252; b = 8'd233;  #10 
a = 8'd252; b = 8'd234;  #10 
a = 8'd252; b = 8'd235;  #10 
a = 8'd252; b = 8'd236;  #10 
a = 8'd252; b = 8'd237;  #10 
a = 8'd252; b = 8'd238;  #10 
a = 8'd252; b = 8'd239;  #10 
a = 8'd252; b = 8'd240;  #10 
a = 8'd252; b = 8'd241;  #10 
a = 8'd252; b = 8'd242;  #10 
a = 8'd252; b = 8'd243;  #10 
a = 8'd252; b = 8'd244;  #10 
a = 8'd252; b = 8'd245;  #10 
a = 8'd252; b = 8'd246;  #10 
a = 8'd252; b = 8'd247;  #10 
a = 8'd252; b = 8'd248;  #10 
a = 8'd252; b = 8'd249;  #10 
a = 8'd252; b = 8'd250;  #10 
a = 8'd252; b = 8'd251;  #10 
a = 8'd252; b = 8'd252;  #10 
a = 8'd252; b = 8'd253;  #10 
a = 8'd252; b = 8'd254;  #10 
a = 8'd252; b = 8'd255;  #10 
a = 8'd253; b = 8'd0;  #10 
a = 8'd253; b = 8'd1;  #10 
a = 8'd253; b = 8'd2;  #10 
a = 8'd253; b = 8'd3;  #10 
a = 8'd253; b = 8'd4;  #10 
a = 8'd253; b = 8'd5;  #10 
a = 8'd253; b = 8'd6;  #10 
a = 8'd253; b = 8'd7;  #10 
a = 8'd253; b = 8'd8;  #10 
a = 8'd253; b = 8'd9;  #10 
a = 8'd253; b = 8'd10;  #10 
a = 8'd253; b = 8'd11;  #10 
a = 8'd253; b = 8'd12;  #10 
a = 8'd253; b = 8'd13;  #10 
a = 8'd253; b = 8'd14;  #10 
a = 8'd253; b = 8'd15;  #10 
a = 8'd253; b = 8'd16;  #10 
a = 8'd253; b = 8'd17;  #10 
a = 8'd253; b = 8'd18;  #10 
a = 8'd253; b = 8'd19;  #10 
a = 8'd253; b = 8'd20;  #10 
a = 8'd253; b = 8'd21;  #10 
a = 8'd253; b = 8'd22;  #10 
a = 8'd253; b = 8'd23;  #10 
a = 8'd253; b = 8'd24;  #10 
a = 8'd253; b = 8'd25;  #10 
a = 8'd253; b = 8'd26;  #10 
a = 8'd253; b = 8'd27;  #10 
a = 8'd253; b = 8'd28;  #10 
a = 8'd253; b = 8'd29;  #10 
a = 8'd253; b = 8'd30;  #10 
a = 8'd253; b = 8'd31;  #10 
a = 8'd253; b = 8'd32;  #10 
a = 8'd253; b = 8'd33;  #10 
a = 8'd253; b = 8'd34;  #10 
a = 8'd253; b = 8'd35;  #10 
a = 8'd253; b = 8'd36;  #10 
a = 8'd253; b = 8'd37;  #10 
a = 8'd253; b = 8'd38;  #10 
a = 8'd253; b = 8'd39;  #10 
a = 8'd253; b = 8'd40;  #10 
a = 8'd253; b = 8'd41;  #10 
a = 8'd253; b = 8'd42;  #10 
a = 8'd253; b = 8'd43;  #10 
a = 8'd253; b = 8'd44;  #10 
a = 8'd253; b = 8'd45;  #10 
a = 8'd253; b = 8'd46;  #10 
a = 8'd253; b = 8'd47;  #10 
a = 8'd253; b = 8'd48;  #10 
a = 8'd253; b = 8'd49;  #10 
a = 8'd253; b = 8'd50;  #10 
a = 8'd253; b = 8'd51;  #10 
a = 8'd253; b = 8'd52;  #10 
a = 8'd253; b = 8'd53;  #10 
a = 8'd253; b = 8'd54;  #10 
a = 8'd253; b = 8'd55;  #10 
a = 8'd253; b = 8'd56;  #10 
a = 8'd253; b = 8'd57;  #10 
a = 8'd253; b = 8'd58;  #10 
a = 8'd253; b = 8'd59;  #10 
a = 8'd253; b = 8'd60;  #10 
a = 8'd253; b = 8'd61;  #10 
a = 8'd253; b = 8'd62;  #10 
a = 8'd253; b = 8'd63;  #10 
a = 8'd253; b = 8'd64;  #10 
a = 8'd253; b = 8'd65;  #10 
a = 8'd253; b = 8'd66;  #10 
a = 8'd253; b = 8'd67;  #10 
a = 8'd253; b = 8'd68;  #10 
a = 8'd253; b = 8'd69;  #10 
a = 8'd253; b = 8'd70;  #10 
a = 8'd253; b = 8'd71;  #10 
a = 8'd253; b = 8'd72;  #10 
a = 8'd253; b = 8'd73;  #10 
a = 8'd253; b = 8'd74;  #10 
a = 8'd253; b = 8'd75;  #10 
a = 8'd253; b = 8'd76;  #10 
a = 8'd253; b = 8'd77;  #10 
a = 8'd253; b = 8'd78;  #10 
a = 8'd253; b = 8'd79;  #10 
a = 8'd253; b = 8'd80;  #10 
a = 8'd253; b = 8'd81;  #10 
a = 8'd253; b = 8'd82;  #10 
a = 8'd253; b = 8'd83;  #10 
a = 8'd253; b = 8'd84;  #10 
a = 8'd253; b = 8'd85;  #10 
a = 8'd253; b = 8'd86;  #10 
a = 8'd253; b = 8'd87;  #10 
a = 8'd253; b = 8'd88;  #10 
a = 8'd253; b = 8'd89;  #10 
a = 8'd253; b = 8'd90;  #10 
a = 8'd253; b = 8'd91;  #10 
a = 8'd253; b = 8'd92;  #10 
a = 8'd253; b = 8'd93;  #10 
a = 8'd253; b = 8'd94;  #10 
a = 8'd253; b = 8'd95;  #10 
a = 8'd253; b = 8'd96;  #10 
a = 8'd253; b = 8'd97;  #10 
a = 8'd253; b = 8'd98;  #10 
a = 8'd253; b = 8'd99;  #10 
a = 8'd253; b = 8'd100;  #10 
a = 8'd253; b = 8'd101;  #10 
a = 8'd253; b = 8'd102;  #10 
a = 8'd253; b = 8'd103;  #10 
a = 8'd253; b = 8'd104;  #10 
a = 8'd253; b = 8'd105;  #10 
a = 8'd253; b = 8'd106;  #10 
a = 8'd253; b = 8'd107;  #10 
a = 8'd253; b = 8'd108;  #10 
a = 8'd253; b = 8'd109;  #10 
a = 8'd253; b = 8'd110;  #10 
a = 8'd253; b = 8'd111;  #10 
a = 8'd253; b = 8'd112;  #10 
a = 8'd253; b = 8'd113;  #10 
a = 8'd253; b = 8'd114;  #10 
a = 8'd253; b = 8'd115;  #10 
a = 8'd253; b = 8'd116;  #10 
a = 8'd253; b = 8'd117;  #10 
a = 8'd253; b = 8'd118;  #10 
a = 8'd253; b = 8'd119;  #10 
a = 8'd253; b = 8'd120;  #10 
a = 8'd253; b = 8'd121;  #10 
a = 8'd253; b = 8'd122;  #10 
a = 8'd253; b = 8'd123;  #10 
a = 8'd253; b = 8'd124;  #10 
a = 8'd253; b = 8'd125;  #10 
a = 8'd253; b = 8'd126;  #10 
a = 8'd253; b = 8'd127;  #10 
a = 8'd253; b = 8'd128;  #10 
a = 8'd253; b = 8'd129;  #10 
a = 8'd253; b = 8'd130;  #10 
a = 8'd253; b = 8'd131;  #10 
a = 8'd253; b = 8'd132;  #10 
a = 8'd253; b = 8'd133;  #10 
a = 8'd253; b = 8'd134;  #10 
a = 8'd253; b = 8'd135;  #10 
a = 8'd253; b = 8'd136;  #10 
a = 8'd253; b = 8'd137;  #10 
a = 8'd253; b = 8'd138;  #10 
a = 8'd253; b = 8'd139;  #10 
a = 8'd253; b = 8'd140;  #10 
a = 8'd253; b = 8'd141;  #10 
a = 8'd253; b = 8'd142;  #10 
a = 8'd253; b = 8'd143;  #10 
a = 8'd253; b = 8'd144;  #10 
a = 8'd253; b = 8'd145;  #10 
a = 8'd253; b = 8'd146;  #10 
a = 8'd253; b = 8'd147;  #10 
a = 8'd253; b = 8'd148;  #10 
a = 8'd253; b = 8'd149;  #10 
a = 8'd253; b = 8'd150;  #10 
a = 8'd253; b = 8'd151;  #10 
a = 8'd253; b = 8'd152;  #10 
a = 8'd253; b = 8'd153;  #10 
a = 8'd253; b = 8'd154;  #10 
a = 8'd253; b = 8'd155;  #10 
a = 8'd253; b = 8'd156;  #10 
a = 8'd253; b = 8'd157;  #10 
a = 8'd253; b = 8'd158;  #10 
a = 8'd253; b = 8'd159;  #10 
a = 8'd253; b = 8'd160;  #10 
a = 8'd253; b = 8'd161;  #10 
a = 8'd253; b = 8'd162;  #10 
a = 8'd253; b = 8'd163;  #10 
a = 8'd253; b = 8'd164;  #10 
a = 8'd253; b = 8'd165;  #10 
a = 8'd253; b = 8'd166;  #10 
a = 8'd253; b = 8'd167;  #10 
a = 8'd253; b = 8'd168;  #10 
a = 8'd253; b = 8'd169;  #10 
a = 8'd253; b = 8'd170;  #10 
a = 8'd253; b = 8'd171;  #10 
a = 8'd253; b = 8'd172;  #10 
a = 8'd253; b = 8'd173;  #10 
a = 8'd253; b = 8'd174;  #10 
a = 8'd253; b = 8'd175;  #10 
a = 8'd253; b = 8'd176;  #10 
a = 8'd253; b = 8'd177;  #10 
a = 8'd253; b = 8'd178;  #10 
a = 8'd253; b = 8'd179;  #10 
a = 8'd253; b = 8'd180;  #10 
a = 8'd253; b = 8'd181;  #10 
a = 8'd253; b = 8'd182;  #10 
a = 8'd253; b = 8'd183;  #10 
a = 8'd253; b = 8'd184;  #10 
a = 8'd253; b = 8'd185;  #10 
a = 8'd253; b = 8'd186;  #10 
a = 8'd253; b = 8'd187;  #10 
a = 8'd253; b = 8'd188;  #10 
a = 8'd253; b = 8'd189;  #10 
a = 8'd253; b = 8'd190;  #10 
a = 8'd253; b = 8'd191;  #10 
a = 8'd253; b = 8'd192;  #10 
a = 8'd253; b = 8'd193;  #10 
a = 8'd253; b = 8'd194;  #10 
a = 8'd253; b = 8'd195;  #10 
a = 8'd253; b = 8'd196;  #10 
a = 8'd253; b = 8'd197;  #10 
a = 8'd253; b = 8'd198;  #10 
a = 8'd253; b = 8'd199;  #10 
a = 8'd253; b = 8'd200;  #10 
a = 8'd253; b = 8'd201;  #10 
a = 8'd253; b = 8'd202;  #10 
a = 8'd253; b = 8'd203;  #10 
a = 8'd253; b = 8'd204;  #10 
a = 8'd253; b = 8'd205;  #10 
a = 8'd253; b = 8'd206;  #10 
a = 8'd253; b = 8'd207;  #10 
a = 8'd253; b = 8'd208;  #10 
a = 8'd253; b = 8'd209;  #10 
a = 8'd253; b = 8'd210;  #10 
a = 8'd253; b = 8'd211;  #10 
a = 8'd253; b = 8'd212;  #10 
a = 8'd253; b = 8'd213;  #10 
a = 8'd253; b = 8'd214;  #10 
a = 8'd253; b = 8'd215;  #10 
a = 8'd253; b = 8'd216;  #10 
a = 8'd253; b = 8'd217;  #10 
a = 8'd253; b = 8'd218;  #10 
a = 8'd253; b = 8'd219;  #10 
a = 8'd253; b = 8'd220;  #10 
a = 8'd253; b = 8'd221;  #10 
a = 8'd253; b = 8'd222;  #10 
a = 8'd253; b = 8'd223;  #10 
a = 8'd253; b = 8'd224;  #10 
a = 8'd253; b = 8'd225;  #10 
a = 8'd253; b = 8'd226;  #10 
a = 8'd253; b = 8'd227;  #10 
a = 8'd253; b = 8'd228;  #10 
a = 8'd253; b = 8'd229;  #10 
a = 8'd253; b = 8'd230;  #10 
a = 8'd253; b = 8'd231;  #10 
a = 8'd253; b = 8'd232;  #10 
a = 8'd253; b = 8'd233;  #10 
a = 8'd253; b = 8'd234;  #10 
a = 8'd253; b = 8'd235;  #10 
a = 8'd253; b = 8'd236;  #10 
a = 8'd253; b = 8'd237;  #10 
a = 8'd253; b = 8'd238;  #10 
a = 8'd253; b = 8'd239;  #10 
a = 8'd253; b = 8'd240;  #10 
a = 8'd253; b = 8'd241;  #10 
a = 8'd253; b = 8'd242;  #10 
a = 8'd253; b = 8'd243;  #10 
a = 8'd253; b = 8'd244;  #10 
a = 8'd253; b = 8'd245;  #10 
a = 8'd253; b = 8'd246;  #10 
a = 8'd253; b = 8'd247;  #10 
a = 8'd253; b = 8'd248;  #10 
a = 8'd253; b = 8'd249;  #10 
a = 8'd253; b = 8'd250;  #10 
a = 8'd253; b = 8'd251;  #10 
a = 8'd253; b = 8'd252;  #10 
a = 8'd253; b = 8'd253;  #10 
a = 8'd253; b = 8'd254;  #10 
a = 8'd253; b = 8'd255;  #10 
a = 8'd254; b = 8'd0;  #10 
a = 8'd254; b = 8'd1;  #10 
a = 8'd254; b = 8'd2;  #10 
a = 8'd254; b = 8'd3;  #10 
a = 8'd254; b = 8'd4;  #10 
a = 8'd254; b = 8'd5;  #10 
a = 8'd254; b = 8'd6;  #10 
a = 8'd254; b = 8'd7;  #10 
a = 8'd254; b = 8'd8;  #10 
a = 8'd254; b = 8'd9;  #10 
a = 8'd254; b = 8'd10;  #10 
a = 8'd254; b = 8'd11;  #10 
a = 8'd254; b = 8'd12;  #10 
a = 8'd254; b = 8'd13;  #10 
a = 8'd254; b = 8'd14;  #10 
a = 8'd254; b = 8'd15;  #10 
a = 8'd254; b = 8'd16;  #10 
a = 8'd254; b = 8'd17;  #10 
a = 8'd254; b = 8'd18;  #10 
a = 8'd254; b = 8'd19;  #10 
a = 8'd254; b = 8'd20;  #10 
a = 8'd254; b = 8'd21;  #10 
a = 8'd254; b = 8'd22;  #10 
a = 8'd254; b = 8'd23;  #10 
a = 8'd254; b = 8'd24;  #10 
a = 8'd254; b = 8'd25;  #10 
a = 8'd254; b = 8'd26;  #10 
a = 8'd254; b = 8'd27;  #10 
a = 8'd254; b = 8'd28;  #10 
a = 8'd254; b = 8'd29;  #10 
a = 8'd254; b = 8'd30;  #10 
a = 8'd254; b = 8'd31;  #10 
a = 8'd254; b = 8'd32;  #10 
a = 8'd254; b = 8'd33;  #10 
a = 8'd254; b = 8'd34;  #10 
a = 8'd254; b = 8'd35;  #10 
a = 8'd254; b = 8'd36;  #10 
a = 8'd254; b = 8'd37;  #10 
a = 8'd254; b = 8'd38;  #10 
a = 8'd254; b = 8'd39;  #10 
a = 8'd254; b = 8'd40;  #10 
a = 8'd254; b = 8'd41;  #10 
a = 8'd254; b = 8'd42;  #10 
a = 8'd254; b = 8'd43;  #10 
a = 8'd254; b = 8'd44;  #10 
a = 8'd254; b = 8'd45;  #10 
a = 8'd254; b = 8'd46;  #10 
a = 8'd254; b = 8'd47;  #10 
a = 8'd254; b = 8'd48;  #10 
a = 8'd254; b = 8'd49;  #10 
a = 8'd254; b = 8'd50;  #10 
a = 8'd254; b = 8'd51;  #10 
a = 8'd254; b = 8'd52;  #10 
a = 8'd254; b = 8'd53;  #10 
a = 8'd254; b = 8'd54;  #10 
a = 8'd254; b = 8'd55;  #10 
a = 8'd254; b = 8'd56;  #10 
a = 8'd254; b = 8'd57;  #10 
a = 8'd254; b = 8'd58;  #10 
a = 8'd254; b = 8'd59;  #10 
a = 8'd254; b = 8'd60;  #10 
a = 8'd254; b = 8'd61;  #10 
a = 8'd254; b = 8'd62;  #10 
a = 8'd254; b = 8'd63;  #10 
a = 8'd254; b = 8'd64;  #10 
a = 8'd254; b = 8'd65;  #10 
a = 8'd254; b = 8'd66;  #10 
a = 8'd254; b = 8'd67;  #10 
a = 8'd254; b = 8'd68;  #10 
a = 8'd254; b = 8'd69;  #10 
a = 8'd254; b = 8'd70;  #10 
a = 8'd254; b = 8'd71;  #10 
a = 8'd254; b = 8'd72;  #10 
a = 8'd254; b = 8'd73;  #10 
a = 8'd254; b = 8'd74;  #10 
a = 8'd254; b = 8'd75;  #10 
a = 8'd254; b = 8'd76;  #10 
a = 8'd254; b = 8'd77;  #10 
a = 8'd254; b = 8'd78;  #10 
a = 8'd254; b = 8'd79;  #10 
a = 8'd254; b = 8'd80;  #10 
a = 8'd254; b = 8'd81;  #10 
a = 8'd254; b = 8'd82;  #10 
a = 8'd254; b = 8'd83;  #10 
a = 8'd254; b = 8'd84;  #10 
a = 8'd254; b = 8'd85;  #10 
a = 8'd254; b = 8'd86;  #10 
a = 8'd254; b = 8'd87;  #10 
a = 8'd254; b = 8'd88;  #10 
a = 8'd254; b = 8'd89;  #10 
a = 8'd254; b = 8'd90;  #10 
a = 8'd254; b = 8'd91;  #10 
a = 8'd254; b = 8'd92;  #10 
a = 8'd254; b = 8'd93;  #10 
a = 8'd254; b = 8'd94;  #10 
a = 8'd254; b = 8'd95;  #10 
a = 8'd254; b = 8'd96;  #10 
a = 8'd254; b = 8'd97;  #10 
a = 8'd254; b = 8'd98;  #10 
a = 8'd254; b = 8'd99;  #10 
a = 8'd254; b = 8'd100;  #10 
a = 8'd254; b = 8'd101;  #10 
a = 8'd254; b = 8'd102;  #10 
a = 8'd254; b = 8'd103;  #10 
a = 8'd254; b = 8'd104;  #10 
a = 8'd254; b = 8'd105;  #10 
a = 8'd254; b = 8'd106;  #10 
a = 8'd254; b = 8'd107;  #10 
a = 8'd254; b = 8'd108;  #10 
a = 8'd254; b = 8'd109;  #10 
a = 8'd254; b = 8'd110;  #10 
a = 8'd254; b = 8'd111;  #10 
a = 8'd254; b = 8'd112;  #10 
a = 8'd254; b = 8'd113;  #10 
a = 8'd254; b = 8'd114;  #10 
a = 8'd254; b = 8'd115;  #10 
a = 8'd254; b = 8'd116;  #10 
a = 8'd254; b = 8'd117;  #10 
a = 8'd254; b = 8'd118;  #10 
a = 8'd254; b = 8'd119;  #10 
a = 8'd254; b = 8'd120;  #10 
a = 8'd254; b = 8'd121;  #10 
a = 8'd254; b = 8'd122;  #10 
a = 8'd254; b = 8'd123;  #10 
a = 8'd254; b = 8'd124;  #10 
a = 8'd254; b = 8'd125;  #10 
a = 8'd254; b = 8'd126;  #10 
a = 8'd254; b = 8'd127;  #10 
a = 8'd254; b = 8'd128;  #10 
a = 8'd254; b = 8'd129;  #10 
a = 8'd254; b = 8'd130;  #10 
a = 8'd254; b = 8'd131;  #10 
a = 8'd254; b = 8'd132;  #10 
a = 8'd254; b = 8'd133;  #10 
a = 8'd254; b = 8'd134;  #10 
a = 8'd254; b = 8'd135;  #10 
a = 8'd254; b = 8'd136;  #10 
a = 8'd254; b = 8'd137;  #10 
a = 8'd254; b = 8'd138;  #10 
a = 8'd254; b = 8'd139;  #10 
a = 8'd254; b = 8'd140;  #10 
a = 8'd254; b = 8'd141;  #10 
a = 8'd254; b = 8'd142;  #10 
a = 8'd254; b = 8'd143;  #10 
a = 8'd254; b = 8'd144;  #10 
a = 8'd254; b = 8'd145;  #10 
a = 8'd254; b = 8'd146;  #10 
a = 8'd254; b = 8'd147;  #10 
a = 8'd254; b = 8'd148;  #10 
a = 8'd254; b = 8'd149;  #10 
a = 8'd254; b = 8'd150;  #10 
a = 8'd254; b = 8'd151;  #10 
a = 8'd254; b = 8'd152;  #10 
a = 8'd254; b = 8'd153;  #10 
a = 8'd254; b = 8'd154;  #10 
a = 8'd254; b = 8'd155;  #10 
a = 8'd254; b = 8'd156;  #10 
a = 8'd254; b = 8'd157;  #10 
a = 8'd254; b = 8'd158;  #10 
a = 8'd254; b = 8'd159;  #10 
a = 8'd254; b = 8'd160;  #10 
a = 8'd254; b = 8'd161;  #10 
a = 8'd254; b = 8'd162;  #10 
a = 8'd254; b = 8'd163;  #10 
a = 8'd254; b = 8'd164;  #10 
a = 8'd254; b = 8'd165;  #10 
a = 8'd254; b = 8'd166;  #10 
a = 8'd254; b = 8'd167;  #10 
a = 8'd254; b = 8'd168;  #10 
a = 8'd254; b = 8'd169;  #10 
a = 8'd254; b = 8'd170;  #10 
a = 8'd254; b = 8'd171;  #10 
a = 8'd254; b = 8'd172;  #10 
a = 8'd254; b = 8'd173;  #10 
a = 8'd254; b = 8'd174;  #10 
a = 8'd254; b = 8'd175;  #10 
a = 8'd254; b = 8'd176;  #10 
a = 8'd254; b = 8'd177;  #10 
a = 8'd254; b = 8'd178;  #10 
a = 8'd254; b = 8'd179;  #10 
a = 8'd254; b = 8'd180;  #10 
a = 8'd254; b = 8'd181;  #10 
a = 8'd254; b = 8'd182;  #10 
a = 8'd254; b = 8'd183;  #10 
a = 8'd254; b = 8'd184;  #10 
a = 8'd254; b = 8'd185;  #10 
a = 8'd254; b = 8'd186;  #10 
a = 8'd254; b = 8'd187;  #10 
a = 8'd254; b = 8'd188;  #10 
a = 8'd254; b = 8'd189;  #10 
a = 8'd254; b = 8'd190;  #10 
a = 8'd254; b = 8'd191;  #10 
a = 8'd254; b = 8'd192;  #10 
a = 8'd254; b = 8'd193;  #10 
a = 8'd254; b = 8'd194;  #10 
a = 8'd254; b = 8'd195;  #10 
a = 8'd254; b = 8'd196;  #10 
a = 8'd254; b = 8'd197;  #10 
a = 8'd254; b = 8'd198;  #10 
a = 8'd254; b = 8'd199;  #10 
a = 8'd254; b = 8'd200;  #10 
a = 8'd254; b = 8'd201;  #10 
a = 8'd254; b = 8'd202;  #10 
a = 8'd254; b = 8'd203;  #10 
a = 8'd254; b = 8'd204;  #10 
a = 8'd254; b = 8'd205;  #10 
a = 8'd254; b = 8'd206;  #10 
a = 8'd254; b = 8'd207;  #10 
a = 8'd254; b = 8'd208;  #10 
a = 8'd254; b = 8'd209;  #10 
a = 8'd254; b = 8'd210;  #10 
a = 8'd254; b = 8'd211;  #10 
a = 8'd254; b = 8'd212;  #10 
a = 8'd254; b = 8'd213;  #10 
a = 8'd254; b = 8'd214;  #10 
a = 8'd254; b = 8'd215;  #10 
a = 8'd254; b = 8'd216;  #10 
a = 8'd254; b = 8'd217;  #10 
a = 8'd254; b = 8'd218;  #10 
a = 8'd254; b = 8'd219;  #10 
a = 8'd254; b = 8'd220;  #10 
a = 8'd254; b = 8'd221;  #10 
a = 8'd254; b = 8'd222;  #10 
a = 8'd254; b = 8'd223;  #10 
a = 8'd254; b = 8'd224;  #10 
a = 8'd254; b = 8'd225;  #10 
a = 8'd254; b = 8'd226;  #10 
a = 8'd254; b = 8'd227;  #10 
a = 8'd254; b = 8'd228;  #10 
a = 8'd254; b = 8'd229;  #10 
a = 8'd254; b = 8'd230;  #10 
a = 8'd254; b = 8'd231;  #10 
a = 8'd254; b = 8'd232;  #10 
a = 8'd254; b = 8'd233;  #10 
a = 8'd254; b = 8'd234;  #10 
a = 8'd254; b = 8'd235;  #10 
a = 8'd254; b = 8'd236;  #10 
a = 8'd254; b = 8'd237;  #10 
a = 8'd254; b = 8'd238;  #10 
a = 8'd254; b = 8'd239;  #10 
a = 8'd254; b = 8'd240;  #10 
a = 8'd254; b = 8'd241;  #10 
a = 8'd254; b = 8'd242;  #10 
a = 8'd254; b = 8'd243;  #10 
a = 8'd254; b = 8'd244;  #10 
a = 8'd254; b = 8'd245;  #10 
a = 8'd254; b = 8'd246;  #10 
a = 8'd254; b = 8'd247;  #10 
a = 8'd254; b = 8'd248;  #10 
a = 8'd254; b = 8'd249;  #10 
a = 8'd254; b = 8'd250;  #10 
a = 8'd254; b = 8'd251;  #10 
a = 8'd254; b = 8'd252;  #10 
a = 8'd254; b = 8'd253;  #10 
a = 8'd254; b = 8'd254;  #10 
a = 8'd254; b = 8'd255;  #10 
a = 8'd255; b = 8'd0;  #10 
a = 8'd255; b = 8'd1;  #10 
a = 8'd255; b = 8'd2;  #10 
a = 8'd255; b = 8'd3;  #10 
a = 8'd255; b = 8'd4;  #10 
a = 8'd255; b = 8'd5;  #10 
a = 8'd255; b = 8'd6;  #10 
a = 8'd255; b = 8'd7;  #10 
a = 8'd255; b = 8'd8;  #10 
a = 8'd255; b = 8'd9;  #10 
a = 8'd255; b = 8'd10;  #10 
a = 8'd255; b = 8'd11;  #10 
a = 8'd255; b = 8'd12;  #10 
a = 8'd255; b = 8'd13;  #10 
a = 8'd255; b = 8'd14;  #10 
a = 8'd255; b = 8'd15;  #10 
a = 8'd255; b = 8'd16;  #10 
a = 8'd255; b = 8'd17;  #10 
a = 8'd255; b = 8'd18;  #10 
a = 8'd255; b = 8'd19;  #10 
a = 8'd255; b = 8'd20;  #10 
a = 8'd255; b = 8'd21;  #10 
a = 8'd255; b = 8'd22;  #10 
a = 8'd255; b = 8'd23;  #10 
a = 8'd255; b = 8'd24;  #10 
a = 8'd255; b = 8'd25;  #10 
a = 8'd255; b = 8'd26;  #10 
a = 8'd255; b = 8'd27;  #10 
a = 8'd255; b = 8'd28;  #10 
a = 8'd255; b = 8'd29;  #10 
a = 8'd255; b = 8'd30;  #10 
a = 8'd255; b = 8'd31;  #10 
a = 8'd255; b = 8'd32;  #10 
a = 8'd255; b = 8'd33;  #10 
a = 8'd255; b = 8'd34;  #10 
a = 8'd255; b = 8'd35;  #10 
a = 8'd255; b = 8'd36;  #10 
a = 8'd255; b = 8'd37;  #10 
a = 8'd255; b = 8'd38;  #10 
a = 8'd255; b = 8'd39;  #10 
a = 8'd255; b = 8'd40;  #10 
a = 8'd255; b = 8'd41;  #10 
a = 8'd255; b = 8'd42;  #10 
a = 8'd255; b = 8'd43;  #10 
a = 8'd255; b = 8'd44;  #10 
a = 8'd255; b = 8'd45;  #10 
a = 8'd255; b = 8'd46;  #10 
a = 8'd255; b = 8'd47;  #10 
a = 8'd255; b = 8'd48;  #10 
a = 8'd255; b = 8'd49;  #10 
a = 8'd255; b = 8'd50;  #10 
a = 8'd255; b = 8'd51;  #10 
a = 8'd255; b = 8'd52;  #10 
a = 8'd255; b = 8'd53;  #10 
a = 8'd255; b = 8'd54;  #10 
a = 8'd255; b = 8'd55;  #10 
a = 8'd255; b = 8'd56;  #10 
a = 8'd255; b = 8'd57;  #10 
a = 8'd255; b = 8'd58;  #10 
a = 8'd255; b = 8'd59;  #10 
a = 8'd255; b = 8'd60;  #10 
a = 8'd255; b = 8'd61;  #10 
a = 8'd255; b = 8'd62;  #10 
a = 8'd255; b = 8'd63;  #10 
a = 8'd255; b = 8'd64;  #10 
a = 8'd255; b = 8'd65;  #10 
a = 8'd255; b = 8'd66;  #10 
a = 8'd255; b = 8'd67;  #10 
a = 8'd255; b = 8'd68;  #10 
a = 8'd255; b = 8'd69;  #10 
a = 8'd255; b = 8'd70;  #10 
a = 8'd255; b = 8'd71;  #10 
a = 8'd255; b = 8'd72;  #10 
a = 8'd255; b = 8'd73;  #10 
a = 8'd255; b = 8'd74;  #10 
a = 8'd255; b = 8'd75;  #10 
a = 8'd255; b = 8'd76;  #10 
a = 8'd255; b = 8'd77;  #10 
a = 8'd255; b = 8'd78;  #10 
a = 8'd255; b = 8'd79;  #10 
a = 8'd255; b = 8'd80;  #10 
a = 8'd255; b = 8'd81;  #10 
a = 8'd255; b = 8'd82;  #10 
a = 8'd255; b = 8'd83;  #10 
a = 8'd255; b = 8'd84;  #10 
a = 8'd255; b = 8'd85;  #10 
a = 8'd255; b = 8'd86;  #10 
a = 8'd255; b = 8'd87;  #10 
a = 8'd255; b = 8'd88;  #10 
a = 8'd255; b = 8'd89;  #10 
a = 8'd255; b = 8'd90;  #10 
a = 8'd255; b = 8'd91;  #10 
a = 8'd255; b = 8'd92;  #10 
a = 8'd255; b = 8'd93;  #10 
a = 8'd255; b = 8'd94;  #10 
a = 8'd255; b = 8'd95;  #10 
a = 8'd255; b = 8'd96;  #10 
a = 8'd255; b = 8'd97;  #10 
a = 8'd255; b = 8'd98;  #10 
a = 8'd255; b = 8'd99;  #10 
a = 8'd255; b = 8'd100;  #10 
a = 8'd255; b = 8'd101;  #10 
a = 8'd255; b = 8'd102;  #10 
a = 8'd255; b = 8'd103;  #10 
a = 8'd255; b = 8'd104;  #10 
a = 8'd255; b = 8'd105;  #10 
a = 8'd255; b = 8'd106;  #10 
a = 8'd255; b = 8'd107;  #10 
a = 8'd255; b = 8'd108;  #10 
a = 8'd255; b = 8'd109;  #10 
a = 8'd255; b = 8'd110;  #10 
a = 8'd255; b = 8'd111;  #10 
a = 8'd255; b = 8'd112;  #10 
a = 8'd255; b = 8'd113;  #10 
a = 8'd255; b = 8'd114;  #10 
a = 8'd255; b = 8'd115;  #10 
a = 8'd255; b = 8'd116;  #10 
a = 8'd255; b = 8'd117;  #10 
a = 8'd255; b = 8'd118;  #10 
a = 8'd255; b = 8'd119;  #10 
a = 8'd255; b = 8'd120;  #10 
a = 8'd255; b = 8'd121;  #10 
a = 8'd255; b = 8'd122;  #10 
a = 8'd255; b = 8'd123;  #10 
a = 8'd255; b = 8'd124;  #10 
a = 8'd255; b = 8'd125;  #10 
a = 8'd255; b = 8'd126;  #10 
a = 8'd255; b = 8'd127;  #10 
a = 8'd255; b = 8'd128;  #10 
a = 8'd255; b = 8'd129;  #10 
a = 8'd255; b = 8'd130;  #10 
a = 8'd255; b = 8'd131;  #10 
a = 8'd255; b = 8'd132;  #10 
a = 8'd255; b = 8'd133;  #10 
a = 8'd255; b = 8'd134;  #10 
a = 8'd255; b = 8'd135;  #10 
a = 8'd255; b = 8'd136;  #10 
a = 8'd255; b = 8'd137;  #10 
a = 8'd255; b = 8'd138;  #10 
a = 8'd255; b = 8'd139;  #10 
a = 8'd255; b = 8'd140;  #10 
a = 8'd255; b = 8'd141;  #10 
a = 8'd255; b = 8'd142;  #10 
a = 8'd255; b = 8'd143;  #10 
a = 8'd255; b = 8'd144;  #10 
a = 8'd255; b = 8'd145;  #10 
a = 8'd255; b = 8'd146;  #10 
a = 8'd255; b = 8'd147;  #10 
a = 8'd255; b = 8'd148;  #10 
a = 8'd255; b = 8'd149;  #10 
a = 8'd255; b = 8'd150;  #10 
a = 8'd255; b = 8'd151;  #10 
a = 8'd255; b = 8'd152;  #10 
a = 8'd255; b = 8'd153;  #10 
a = 8'd255; b = 8'd154;  #10 
a = 8'd255; b = 8'd155;  #10 
a = 8'd255; b = 8'd156;  #10 
a = 8'd255; b = 8'd157;  #10 
a = 8'd255; b = 8'd158;  #10 
a = 8'd255; b = 8'd159;  #10 
a = 8'd255; b = 8'd160;  #10 
a = 8'd255; b = 8'd161;  #10 
a = 8'd255; b = 8'd162;  #10 
a = 8'd255; b = 8'd163;  #10 
a = 8'd255; b = 8'd164;  #10 
a = 8'd255; b = 8'd165;  #10 
a = 8'd255; b = 8'd166;  #10 
a = 8'd255; b = 8'd167;  #10 
a = 8'd255; b = 8'd168;  #10 
a = 8'd255; b = 8'd169;  #10 
a = 8'd255; b = 8'd170;  #10 
a = 8'd255; b = 8'd171;  #10 
a = 8'd255; b = 8'd172;  #10 
a = 8'd255; b = 8'd173;  #10 
a = 8'd255; b = 8'd174;  #10 
a = 8'd255; b = 8'd175;  #10 
a = 8'd255; b = 8'd176;  #10 
a = 8'd255; b = 8'd177;  #10 
a = 8'd255; b = 8'd178;  #10 
a = 8'd255; b = 8'd179;  #10 
a = 8'd255; b = 8'd180;  #10 
a = 8'd255; b = 8'd181;  #10 
a = 8'd255; b = 8'd182;  #10 
a = 8'd255; b = 8'd183;  #10 
a = 8'd255; b = 8'd184;  #10 
a = 8'd255; b = 8'd185;  #10 
a = 8'd255; b = 8'd186;  #10 
a = 8'd255; b = 8'd187;  #10 
a = 8'd255; b = 8'd188;  #10 
a = 8'd255; b = 8'd189;  #10 
a = 8'd255; b = 8'd190;  #10 
a = 8'd255; b = 8'd191;  #10 
a = 8'd255; b = 8'd192;  #10 
a = 8'd255; b = 8'd193;  #10 
a = 8'd255; b = 8'd194;  #10 
a = 8'd255; b = 8'd195;  #10 
a = 8'd255; b = 8'd196;  #10 
a = 8'd255; b = 8'd197;  #10 
a = 8'd255; b = 8'd198;  #10 
a = 8'd255; b = 8'd199;  #10 
a = 8'd255; b = 8'd200;  #10 
a = 8'd255; b = 8'd201;  #10 
a = 8'd255; b = 8'd202;  #10 
a = 8'd255; b = 8'd203;  #10 
a = 8'd255; b = 8'd204;  #10 
a = 8'd255; b = 8'd205;  #10 
a = 8'd255; b = 8'd206;  #10 
a = 8'd255; b = 8'd207;  #10 
a = 8'd255; b = 8'd208;  #10 
a = 8'd255; b = 8'd209;  #10 
a = 8'd255; b = 8'd210;  #10 
a = 8'd255; b = 8'd211;  #10 
a = 8'd255; b = 8'd212;  #10 
a = 8'd255; b = 8'd213;  #10 
a = 8'd255; b = 8'd214;  #10 
a = 8'd255; b = 8'd215;  #10 
a = 8'd255; b = 8'd216;  #10 
a = 8'd255; b = 8'd217;  #10 
a = 8'd255; b = 8'd218;  #10 
a = 8'd255; b = 8'd219;  #10 
a = 8'd255; b = 8'd220;  #10 
a = 8'd255; b = 8'd221;  #10 
a = 8'd255; b = 8'd222;  #10 
a = 8'd255; b = 8'd223;  #10 
a = 8'd255; b = 8'd224;  #10 
a = 8'd255; b = 8'd225;  #10 
a = 8'd255; b = 8'd226;  #10 
a = 8'd255; b = 8'd227;  #10 
a = 8'd255; b = 8'd228;  #10 
a = 8'd255; b = 8'd229;  #10 
a = 8'd255; b = 8'd230;  #10 
a = 8'd255; b = 8'd231;  #10 
a = 8'd255; b = 8'd232;  #10 
a = 8'd255; b = 8'd233;  #10 
a = 8'd255; b = 8'd234;  #10 
a = 8'd255; b = 8'd235;  #10 
a = 8'd255; b = 8'd236;  #10 
a = 8'd255; b = 8'd237;  #10 
a = 8'd255; b = 8'd238;  #10 
a = 8'd255; b = 8'd239;  #10 
a = 8'd255; b = 8'd240;  #10 
a = 8'd255; b = 8'd241;  #10 
a = 8'd255; b = 8'd242;  #10 
a = 8'd255; b = 8'd243;  #10 
a = 8'd255; b = 8'd244;  #10 
a = 8'd255; b = 8'd245;  #10 
a = 8'd255; b = 8'd246;  #10 
a = 8'd255; b = 8'd247;  #10 
a = 8'd255; b = 8'd248;  #10 
a = 8'd255; b = 8'd249;  #10 
a = 8'd255; b = 8'd250;  #10 
a = 8'd255; b = 8'd251;  #10 
a = 8'd255; b = 8'd252;  #10 
a = 8'd255; b = 8'd253;  #10 
a = 8'd255; b = 8'd254;  #10 
a = 8'd255; b = 8'd255;  #10 

;end


 initial 

 begin 
$monitor("  a,b,product  %d , %d , %d , ",a,b,product) ;
end

endmodule