//check this
// input t1;
// input t1 ;
module not;
