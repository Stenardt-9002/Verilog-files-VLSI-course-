module assing1mod (inp1,ouy1);
input [10:0]inp1;
output [10:0]ouy1;

  assign ouy1 = inp1;

endmodule // assing1mod
